
module CONV_DW01_add_0 ( A, B, CI, SUM, CO );
  input [43:0] A;
  input [43:0] B;
  output [43:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19;
  wire   [43:1] carry;
  assign SUM[19] = A[19];
  assign SUM[18] = A[18];
  assign SUM[17] = A[17];
  assign SUM[16] = A[16];
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  XOR2X1 U1 ( .A(A[40]), .B(n15), .Y(SUM[40]) );
  XOR2X1 U2 ( .A(A[42]), .B(n13), .Y(SUM[42]) );
  XOR2X1 U3 ( .A(A[41]), .B(n14), .Y(SUM[41]) );
  XOR2X1 U4 ( .A(A[39]), .B(n16), .Y(SUM[39]) );
  XOR2X1 U5 ( .A(A[34]), .B(n5), .Y(SUM[34]) );
  XOR2X1 U6 ( .A(A[31]), .B(n8), .Y(SUM[31]) );
  XOR2X1 U7 ( .A(A[30]), .B(n9), .Y(SUM[30]) );
  XOR2X1 U8 ( .A(A[29]), .B(carry[29]), .Y(SUM[29]) );
  XNOR2X1 U9 ( .A(A[28]), .B(n2), .Y(SUM[28]) );
  XOR2X1 U10 ( .A(A[23]), .B(n11), .Y(SUM[23]) );
  XOR2X1 U11 ( .A(A[38]), .B(n17), .Y(SUM[38]) );
  XOR2X1 U12 ( .A(A[37]), .B(n18), .Y(SUM[37]) );
  XOR2X1 U13 ( .A(A[36]), .B(n12), .Y(SUM[36]) );
  XOR2X1 U14 ( .A(A[35]), .B(n4), .Y(SUM[35]) );
  XOR2X1 U15 ( .A(A[33]), .B(n6), .Y(SUM[33]) );
  XOR2X1 U16 ( .A(A[27]), .B(n10), .Y(SUM[27]) );
  XOR2X1 U17 ( .A(A[26]), .B(carry[26]), .Y(SUM[26]) );
  XNOR2X1 U18 ( .A(A[25]), .B(carry[25]), .Y(SUM[25]) );
  XNOR2X1 U19 ( .A(A[24]), .B(n3), .Y(SUM[24]) );
  XOR2X1 U20 ( .A(A[32]), .B(n7), .Y(SUM[32]) );
  XOR2X1 U21 ( .A(A[22]), .B(n1), .Y(SUM[22]) );
  XOR2X1 U22 ( .A(A[21]), .B(A[20]), .Y(SUM[21]) );
  CLKINVX1 U23 ( .A(A[20]), .Y(SUM[20]) );
  XNOR2X1 U24 ( .A(A[43]), .B(n19), .Y(SUM[43]) );
  NAND2X1 U25 ( .A(A[42]), .B(n13), .Y(n19) );
  OR2X1 U26 ( .A(A[24]), .B(n3), .Y(carry[25]) );
  OR2X1 U27 ( .A(A[28]), .B(n2), .Y(carry[29]) );
  OR2X1 U28 ( .A(A[25]), .B(carry[25]), .Y(carry[26]) );
  AND2X2 U29 ( .A(A[21]), .B(A[20]), .Y(n1) );
  AND2X2 U30 ( .A(A[27]), .B(n10), .Y(n2) );
  AND2X2 U31 ( .A(A[23]), .B(n11), .Y(n3) );
  AND2X2 U32 ( .A(A[34]), .B(n5), .Y(n4) );
  AND2X2 U33 ( .A(A[33]), .B(n6), .Y(n5) );
  AND2X2 U34 ( .A(A[32]), .B(n7), .Y(n6) );
  AND2X2 U35 ( .A(A[31]), .B(n8), .Y(n7) );
  AND2X2 U36 ( .A(A[30]), .B(n9), .Y(n8) );
  AND2X2 U37 ( .A(A[29]), .B(carry[29]), .Y(n9) );
  AND2X2 U38 ( .A(A[26]), .B(carry[26]), .Y(n10) );
  AND2X2 U39 ( .A(A[22]), .B(n1), .Y(n11) );
  AND2X2 U40 ( .A(A[35]), .B(n4), .Y(n12) );
  AND2X2 U41 ( .A(A[41]), .B(n14), .Y(n13) );
  AND2X2 U42 ( .A(A[40]), .B(n15), .Y(n14) );
  AND2X2 U43 ( .A(A[39]), .B(n16), .Y(n15) );
  AND2X2 U44 ( .A(A[38]), .B(n17), .Y(n16) );
  AND2X2 U45 ( .A(A[37]), .B(n18), .Y(n17) );
  AND2X2 U46 ( .A(A[36]), .B(n12), .Y(n18) );
endmodule


module CONV_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [19:0] A;
  input [19:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178;

  AOI221X1 U55 ( .A0(A[10]), .A1(n124), .B0(n155), .B1(n156), .C0(n157), .Y(
        n144) );
  OAI222X2 U56 ( .A0(B[12]), .A1(n122), .B0(B[12]), .B1(n150), .C0(n122), .C1(
        n150), .Y(n149) );
  NAND2X4 U57 ( .A(A[11]), .B(n132), .Y(n150) );
  OAI222X1 U58 ( .A0(A[6]), .A1(n165), .B0(n134), .B1(n165), .C0(A[6]), .C1(
        n134), .Y(n164) );
  OAI222X1 U59 ( .A0(B[5]), .A1(n126), .B0(B[5]), .B1(n166), .C0(n126), .C1(
        n166), .Y(n165) );
  OAI222X1 U60 ( .A0(A[13]), .A1(n153), .B0(n153), .B1(n131), .C0(A[13]), .C1(
        n131), .Y(n152) );
  OAI222X4 U61 ( .A0(B[12]), .A1(n122), .B0(B[12]), .B1(n154), .C0(n154), .C1(
        n122), .Y(n153) );
  OAI221X1 U62 ( .A0(B[19]), .A1(n137), .B0(B[19]), .B1(n119), .C0(n138), .Y(
        GE_LT_GT_LE) );
  OAI22X2 U63 ( .A0(n123), .A1(n159), .B0(B[10]), .B1(n159), .Y(n156) );
  OAI21X2 U64 ( .A0(A[9]), .A1(n133), .B0(n160), .Y(n159) );
  OAI22X1 U65 ( .A0(n173), .A1(n127), .B0(B[3]), .B1(n173), .Y(n170) );
  NOR2BX1 U66 ( .AN(B[2]), .B(A[2]), .Y(n173) );
  OAI22X2 U67 ( .A0(B[10]), .A1(n123), .B0(B[10]), .B1(n158), .Y(n157) );
  INVX2 U68 ( .A(n158), .Y(n124) );
  OAI222X4 U69 ( .A0(A[9]), .A1(n175), .B0(n175), .B1(n133), .C0(A[9]), .C1(
        n133), .Y(n158) );
  INVX8 U70 ( .A(A[12]), .Y(n122) );
  OAI21X1 U71 ( .A0(n144), .A1(n145), .B0(n146), .Y(n139) );
  OAI222X1 U72 ( .A0(A[15]), .A1(n147), .B0(n130), .B1(n147), .C0(A[15]), .C1(
        n130), .Y(n146) );
  OAI222XL U73 ( .A0(B[14]), .A1(n121), .B0(B[14]), .B1(n148), .C0(n121), .C1(
        n148), .Y(n147) );
  OAI222XL U74 ( .A0(B[17]), .A1(n120), .B0(B[17]), .B1(n178), .C0(n178), .C1(
        n120), .Y(n177) );
  OAI222X1 U75 ( .A0(A[13]), .A1(n149), .B0(n131), .B1(n149), .C0(A[13]), .C1(
        n131), .Y(n148) );
  CLKINVX1 U76 ( .A(B[13]), .Y(n131) );
  NAND2BXL U77 ( .AN(B[7]), .B(A[7]), .Y(n176) );
  NOR2BXL U78 ( .AN(B[7]), .B(A[7]), .Y(n161) );
  OAI222X4 U79 ( .A0(B[8]), .A1(n125), .B0(B[8]), .B1(n176), .C0(n176), .C1(
        n125), .Y(n175) );
  NAND2BXL U80 ( .AN(B[2]), .B(A[2]), .Y(n172) );
  AOI2BB1XL U81 ( .A0N(n136), .A1N(A[1]), .B0(B[0]), .Y(n174) );
  NAND2BXL U82 ( .AN(B[16]), .B(A[16]), .Y(n178) );
  NOR2BXL U83 ( .AN(B[16]), .B(A[16]), .Y(n143) );
  AOI2BB2X1 U84 ( .B0(n139), .B1(n140), .A0N(n137), .A1N(n119), .Y(n138) );
  CLKINVX1 U85 ( .A(n172), .Y(n128) );
  INVXL U86 ( .A(B[1]), .Y(n136) );
  CLKINVX1 U87 ( .A(A[5]), .Y(n126) );
  CLKINVX1 U88 ( .A(A[8]), .Y(n125) );
  CLKINVX1 U89 ( .A(A[14]), .Y(n121) );
  CLKINVX1 U90 ( .A(A[17]), .Y(n120) );
  CLKINVX1 U91 ( .A(A[3]), .Y(n127) );
  CLKINVX1 U92 ( .A(A[10]), .Y(n123) );
  INVXL U93 ( .A(B[11]), .Y(n132) );
  CLKINVX1 U94 ( .A(A[19]), .Y(n119) );
  INVXL U95 ( .A(B[9]), .Y(n133) );
  INVXL U96 ( .A(B[4]), .Y(n135) );
  INVXL U97 ( .A(B[6]), .Y(n134) );
  INVXL U98 ( .A(B[18]), .Y(n129) );
  INVXL U99 ( .A(B[15]), .Y(n130) );
  OAI22XL U100 ( .A0(n119), .A1(n141), .B0(B[19]), .B1(n141), .Y(n140) );
  OAI21XL U101 ( .A0(A[18]), .A1(n129), .B0(n142), .Y(n141) );
  OAI22XL U102 ( .A0(n143), .A1(n120), .B0(B[17]), .B1(n143), .Y(n142) );
  OAI21XL U103 ( .A0(A[15]), .A1(n130), .B0(n151), .Y(n145) );
  OAI22XL U104 ( .A0(n152), .A1(n121), .B0(B[14]), .B1(n152), .Y(n151) );
  NOR2X1 U105 ( .A(n132), .B(A[11]), .Y(n154) );
  OAI22XL U106 ( .A0(n161), .A1(n125), .B0(B[8]), .B1(n161), .Y(n160) );
  OAI21XL U107 ( .A0(n162), .A1(n163), .B0(n164), .Y(n155) );
  NAND2X1 U108 ( .A(A[4]), .B(n135), .Y(n166) );
  OAI21XL U109 ( .A0(A[6]), .A1(n134), .B0(n167), .Y(n163) );
  OAI22XL U110 ( .A0(n168), .A1(n126), .B0(B[5]), .B1(n168), .Y(n167) );
  NOR2X1 U111 ( .A(n135), .B(A[4]), .Y(n168) );
  AOI221XL U112 ( .A0(A[3]), .A1(n128), .B0(n169), .B1(n170), .C0(n171), .Y(
        n162) );
  OAI22XL U113 ( .A0(B[3]), .A1(n127), .B0(B[3]), .B1(n172), .Y(n171) );
  AO22X1 U114 ( .A0(n174), .A1(A[0]), .B0(A[1]), .B1(n136), .Y(n169) );
  OAI222XL U115 ( .A0(A[18]), .A1(n177), .B0(n177), .B1(n129), .C0(A[18]), 
        .C1(n129), .Y(n137) );
endmodule


module CONV_DW01_inc_0 ( A, SUM );
  input [20:0] A;
  output [20:0] SUM;

  wire   [20:2] carry;

  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR2X1 U1 ( .A(carry[20]), .B(A[20]), .Y(SUM[20]) );
endmodule


module CONV_DW_mult_tc_2 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n3, n6, n7, n9, n11, n12, n13, n15, n16, n17, n18, n19, n21, n22,
         n23, n24, n25, n28, n30, n31, n34, n35, n36, n37, n39, n40, n41, n43,
         n46, n47, n49, n52, n54, n55, n57, n58, n59, n60, n61, n63, n65, n66,
         n67, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n101, n102, n103, n104, n106, n108, n109, n110, n111, n112,
         n113, n115, n116, n117, n118, n120, n122, n123, n124, n125, n126,
         n127, n129, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n152, n153, n154,
         n155, n156, n158, n160, n161, n163, n165, n167, n168, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n183,
         n184, n185, n186, n187, n188, n190, n192, n193, n194, n195, n196,
         n197, n198, n200, n201, n202, n203, n204, n205, n206, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n225, n226, n227, n228, n229, n230, n231, n232, n234, n235, n236,
         n237, n238, n239, n240, n241, n244, n246, n247, n248, n249, n250,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n271, n272, n273, n274,
         n275, n276, n277, n280, n281, n282, n283, n284, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n297, n299, n302, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n324, n326, n327, n328, n330,
         n332, n333, n334, n335, n336, n337, n338, n339, n342, n344, n345,
         n346, n348, n350, n351, n352, n353, n354, n355, n357, n360, n367,
         n369, n371, n372, n373, n375, n376, n377, n378, n381, n382, n389,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         \product[39] , n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197;
  assign product[37] = n101;
  assign product[38] = n101;
  assign product[36] = \product[39] ;
  assign product[39] = \product[39] ;

  BUFX4 U949 ( .A(n812), .Y(n1127) );
  OAI22X2 U950 ( .A0(n915), .A1(n24), .B0(n914), .B1(n22), .Y(n736) );
  BUFX4 U951 ( .A(n807), .Y(n1122) );
  XNOR2X2 U952 ( .A(n988), .B(n31), .Y(n880) );
  OAI22X2 U953 ( .A0(n879), .A1(n36), .B0(n878), .B1(n34), .Y(n701) );
  CLKXOR2X2 U954 ( .A(n314), .B(n89), .Y(product[9]) );
  BUFX4 U955 ( .A(n956), .Y(n1123) );
  NOR2X2 U956 ( .A(n566), .B(n575), .Y(n290) );
  BUFX4 U957 ( .A(n1026), .Y(n34) );
  XNOR2X1 U958 ( .A(n991), .B(n25), .Y(n901) );
  OAI22X1 U959 ( .A0(n946), .A1(n17), .B0(n945), .B1(n15), .Y(n767) );
  OAI22X1 U960 ( .A0(n944), .A1(n15), .B0(n945), .B1(n17), .Y(n766) );
  XNOR2X2 U961 ( .A(a[2]), .B(n13), .Y(n945) );
  OAI22X1 U962 ( .A0(n852), .A1(n46), .B0(n853), .B1(n47), .Y(n677) );
  XNOR2X2 U963 ( .A(n996), .B(n7), .Y(n960) );
  BUFX6 U964 ( .A(a[5]), .Y(n996) );
  BUFX3 U965 ( .A(n641), .Y(n1124) );
  AOI21X2 U966 ( .A0(n258), .A1(n275), .B0(n259), .Y(n257) );
  OAI21X1 U967 ( .A0(n260), .A1(n268), .B0(n261), .Y(n259) );
  CMPR42X2 U968 ( .A(n709), .B(n530), .C(n539), .D(n724), .ICI(n540), .S(n525), 
        .ICO(n523), .CO(n524) );
  OAI22X1 U969 ( .A0(n887), .A1(n35), .B0(n886), .B1(n34), .Y(n709) );
  XNOR2X1 U970 ( .A(n986), .B(n13), .Y(n932) );
  CLKBUFX6 U971 ( .A(a[15]), .Y(n986) );
  XNOR2X2 U972 ( .A(b[16]), .B(b[15]), .Y(n1023) );
  BUFX4 U973 ( .A(b[17]), .Y(n49) );
  OAI22X1 U974 ( .A0(n864), .A1(n41), .B0(n863), .B1(n40), .Y(n687) );
  BUFX6 U975 ( .A(n1015), .Y(n41) );
  XNOR2X1 U976 ( .A(n988), .B(n43), .Y(n844) );
  BUFX6 U977 ( .A(a[13]), .Y(n988) );
  XNOR2X1 U978 ( .A(n989), .B(n37), .Y(n863) );
  CLKBUFX3 U979 ( .A(n692), .Y(n1125) );
  XNOR2X2 U980 ( .A(n992), .B(n49), .Y(n830) );
  OAI22X2 U981 ( .A0(n815), .A1(n57), .B0(n816), .B1(n59), .Y(n644) );
  XNOR2X1 U982 ( .A(b[4]), .B(b[3]), .Y(n1029) );
  CLKBUFX3 U983 ( .A(b[3]), .Y(n7) );
  OAI22X1 U984 ( .A0(n898), .A1(n28), .B0(n899), .B1(n30), .Y(n720) );
  XNOR2X1 U985 ( .A(n988), .B(n25), .Y(n898) );
  OAI22X1 U986 ( .A0(n869), .A1(n39), .B0(n870), .B1(n41), .Y(n693) );
  CLKBUFX3 U987 ( .A(n707), .Y(n1126) );
  OAI22XL U988 ( .A0(n880), .A1(n34), .B0(n881), .B1(n36), .Y(n703) );
  OAI22X1 U989 ( .A0(n882), .A1(n36), .B0(n881), .B1(n34), .Y(n704) );
  CMPR42X1 U990 ( .A(n693), .B(n529), .C(n723), .D(n755), .ICI(n523), .S(n512), 
        .ICO(n510), .CO(n511) );
  OAI22X1 U991 ( .A0(n902), .A1(n30), .B0(n901), .B1(n28), .Y(n723) );
  XNOR2X1 U992 ( .A(n991), .B(n1), .Y(n973) );
  BUFX3 U993 ( .A(n689), .Y(n1128) );
  OAI22X1 U994 ( .A0(n1131), .A1(n47), .B0(n847), .B1(n46), .Y(n672) );
  BUFX4 U995 ( .A(n848), .Y(n1131) );
  OAI22X2 U996 ( .A0(n818), .A1(n57), .B0(n819), .B1(n59), .Y(n646) );
  XNOR2X2 U997 ( .A(a[2]), .B(n55), .Y(n819) );
  NAND2X2 U998 ( .A(n1166), .B(n1167), .Y(product[21]) );
  OAI22X2 U999 ( .A0(n896), .A1(n30), .B0(n895), .B1(n28), .Y(n449) );
  OAI22X2 U1000 ( .A0(n906), .A1(n28), .B0(n907), .B1(n30), .Y(n728) );
  OAI22X2 U1001 ( .A0(n908), .A1(n28), .B0(n909), .B1(n30), .Y(n730) );
  BUFX4 U1002 ( .A(n1027), .Y(n28) );
  BUFX8 U1003 ( .A(n920), .Y(n1129) );
  XNOR2X1 U1004 ( .A(n992), .B(n19), .Y(n920) );
  CMPR42X2 U1005 ( .A(n432), .B(n670), .C(n642), .D(n439), .ICI(n656), .S(n430), .ICO(n428), .CO(n429) );
  OAI22XL U1006 ( .A0(n902), .A1(n28), .B0(n903), .B1(n30), .Y(n724) );
  OAI22XL U1007 ( .A0(n910), .A1(n28), .B0(n911), .B1(n30), .Y(n732) );
  OAI22XL U1008 ( .A0(n900), .A1(n28), .B0(n901), .B1(n30), .Y(n722) );
  OAI22X1 U1009 ( .A0(n905), .A1(n28), .B0(n906), .B1(n30), .Y(n727) );
  OAI22X1 U1010 ( .A0(n907), .A1(n28), .B0(n908), .B1(n1017), .Y(n729) );
  XNOR2X4 U1011 ( .A(n193), .B(n72), .Y(product[26]) );
  BUFX12 U1012 ( .A(a[0]), .Y(n61) );
  CMPR42X2 U1013 ( .A(n624), .B(n754), .C(n648), .D(n516), .ICI(n513), .S(n503), .ICO(n501), .CO(n502) );
  OAI22X1 U1014 ( .A0(n822), .A1(n58), .B0(n60), .B1(n1032), .Y(n624) );
  XNOR2X4 U1015 ( .A(a[1]), .B(n55), .Y(n820) );
  XNOR2X1 U1016 ( .A(n991), .B(n31), .Y(n883) );
  CMPR42X2 U1017 ( .A(n790), .B(n681), .C(n726), .D(n742), .ICI(n562), .S(n549), .ICO(n547), .CO(n548) );
  OAI22X1 U1018 ( .A0(n969), .A1(n6), .B0(n968), .B1(n3), .Y(n790) );
  CMPR42X2 U1019 ( .A(n676), .B(n706), .C(n737), .D(n501), .ICI(n498), .S(n487), .ICO(n485), .CO(n486) );
  OAI22X1 U1020 ( .A0(n851), .A1(n46), .B0(n852), .B1(n47), .Y(n676) );
  XOR2X4 U1021 ( .A(n269), .B(n81), .Y(product[17]) );
  OAI22X1 U1022 ( .A0(n936), .A1(n16), .B0(n937), .B1(n18), .Y(n758) );
  ADDFHX2 U1023 ( .A(n619), .B(n631), .CI(n768), .CO(n616), .S(n617) );
  ADDHX1 U1024 ( .A(n784), .B(n800), .CO(n618), .S(n619) );
  BUFX8 U1025 ( .A(n830), .Y(n1130) );
  NAND2X4 U1026 ( .A(n1173), .B(n1174), .Y(n902) );
  XNOR2X4 U1027 ( .A(n1194), .B(n93), .Y(product[5]) );
  OAI22X1 U1028 ( .A0(n820), .A1(n57), .B0(n821), .B1(n59), .Y(n648) );
  OAI22X1 U1029 ( .A0(n1131), .A1(n46), .B0(n849), .B1(n47), .Y(n673) );
  OAI22X1 U1030 ( .A0(n860), .A1(n41), .B0(n859), .B1(n40), .Y(n417) );
  XNOR2X1 U1031 ( .A(n985), .B(n37), .Y(n859) );
  OAI22X1 U1032 ( .A0(n858), .A1(n46), .B0(n47), .B1(n1183), .Y(n626) );
  OAI22X1 U1033 ( .A0(n833), .A1(n52), .B0(n834), .B1(n1013), .Y(n660) );
  OAI22X1 U1034 ( .A0(n856), .A1(n1024), .B0(n857), .B1(n47), .Y(n681) );
  CMPR42X2 U1035 ( .A(n701), .B(n440), .C(n447), .D(n657), .ICI(n444), .S(n438), .ICO(n436), .CO(n437) );
  OAI22X1 U1036 ( .A0(n946), .A1(n15), .B0(n947), .B1(n17), .Y(n768) );
  XNOR2XL U1037 ( .A(n61), .B(n13), .Y(n947) );
  BUFX8 U1038 ( .A(n247), .Y(n1132) );
  NOR2X2 U1039 ( .A(n252), .B(n249), .Y(n247) );
  XOR2X4 U1040 ( .A(n262), .B(n80), .Y(product[18]) );
  CMPR42X2 U1041 ( .A(n658), .B(n644), .C(n448), .D(n672), .ICI(n458), .S(n446), .ICO(n444), .CO(n445) );
  OAI22X2 U1042 ( .A0(n978), .A1(n3), .B0(n979), .B1(n6), .Y(n800) );
  AO21X2 U1043 ( .A0(n6), .A1(n3), .B0(n967), .Y(n788) );
  OAI22X2 U1044 ( .A0(n980), .A1(n3), .B0(n981), .B1(n6), .Y(n802) );
  OAI22X2 U1045 ( .A0(n982), .A1(n6), .B0(n981), .B1(n3), .Y(n803) );
  BUFX4 U1046 ( .A(n1021), .Y(n6) );
  OAI22X1 U1047 ( .A0(n964), .A1(n9), .B0(n965), .B1(n11), .Y(n786) );
  XNOR2XL U1048 ( .A(n61), .B(n7), .Y(n965) );
  XOR2X4 U1049 ( .A(n322), .B(n90), .Y(product[8]) );
  XNOR2X2 U1050 ( .A(n351), .B(n95), .Y(product[3]) );
  AOI21X2 U1051 ( .A0(n351), .A1(n1142), .B0(n348), .Y(n346) );
  OAI21X1 U1052 ( .A0(n352), .A1(n355), .B0(n353), .Y(n351) );
  NAND2X1 U1053 ( .A(n786), .B(n623), .Y(n350) );
  ADDHX2 U1054 ( .A(n802), .B(n632), .CO(n622), .S(n623) );
  BUFX4 U1055 ( .A(a[11]), .Y(n990) );
  CLKINVX3 U1056 ( .A(n160), .Y(n158) );
  OAI22XL U1057 ( .A0(n900), .A1(n30), .B0(n899), .B1(n28), .Y(n721) );
  XNOR2X1 U1058 ( .A(n990), .B(n43), .Y(n846) );
  OAI22XL U1059 ( .A0(n897), .A1(n30), .B0(n896), .B1(n28), .Y(n718) );
  OAI22X1 U1060 ( .A0(n888), .A1(n34), .B0(n889), .B1(n35), .Y(n711) );
  OAI22X1 U1061 ( .A0(n853), .A1(n46), .B0(n854), .B1(n47), .Y(n678) );
  NAND2X1 U1062 ( .A(n1175), .B(n1176), .Y(n739) );
  OAI22X1 U1063 ( .A0(n840), .A1(n52), .B0(n54), .B1(n1159), .Y(n625) );
  OAI22X1 U1064 ( .A0(n926), .A1(n21), .B0(n927), .B1(n23), .Y(n748) );
  OAI22XL U1065 ( .A0(n856), .A1(n47), .B0(n855), .B1(n1024), .Y(n680) );
  OAI22XL U1066 ( .A0(n838), .A1(n52), .B0(n839), .B1(n1013), .Y(n664) );
  OAI22XL U1067 ( .A0(n951), .A1(n12), .B0(n950), .B1(n9), .Y(n772) );
  CLKINVX1 U1068 ( .A(n122), .Y(n120) );
  CLKINVX1 U1069 ( .A(n165), .Y(n163) );
  INVX3 U1070 ( .A(n293), .Y(n1190) );
  OAI22X1 U1071 ( .A0(n846), .A1(n46), .B0(n847), .B1(n47), .Y(n671) );
  OAI22XL U1072 ( .A0(n898), .A1(n30), .B0(n897), .B1(n28), .Y(n719) );
  NOR2X1 U1073 ( .A(n473), .B(n483), .Y(n238) );
  ADDFXL U1074 ( .A(n683), .B(n417), .CI(n639), .CO(n410), .S(n411) );
  OAI22XL U1075 ( .A0(n954), .A1(n9), .B0(n955), .B1(n12), .Y(n776) );
  OR2X2 U1076 ( .A(n960), .B(n9), .Y(n1195) );
  CLKINVX1 U1077 ( .A(n192), .Y(n190) );
  CMPR42X1 U1078 ( .A(n479), .B(n489), .C(n486), .D(n476), .ICI(n482), .S(n473), .ICO(n471), .CO(n472) );
  CMPR42X1 U1079 ( .A(n467), .B(n459), .C(n464), .D(n456), .ICI(n460), .S(n453), .ICO(n451), .CO(n452) );
  OAI22XL U1080 ( .A0(n904), .A1(n30), .B0(n903), .B1(n28), .Y(n725) );
  ADDFXL U1081 ( .A(n398), .B(n636), .CI(n399), .CO(n395), .S(n396) );
  OAI22XL U1082 ( .A0(n838), .A1(n1013), .B0(n837), .B1(n52), .Y(n663) );
  OAI22XL U1083 ( .A0(n886), .A1(n35), .B0(n885), .B1(n34), .Y(n708) );
  OAI22XL U1084 ( .A0(n934), .A1(n18), .B0(n933), .B1(n16), .Y(n755) );
  OAI22XL U1085 ( .A0(n940), .A1(n17), .B0(n939), .B1(n15), .Y(n761) );
  CMPR42X1 U1086 ( .A(n589), .B(n794), .C(n628), .D(n593), .ICI(n778), .S(n587), .ICO(n585), .CO(n586) );
  OAI22XL U1087 ( .A0(n972), .A1(n3), .B0(n973), .B1(n6), .Y(n794) );
  BUFX4 U1088 ( .A(b[11]), .Y(n31) );
  XOR2X1 U1089 ( .A(b[0]), .B(b[1]), .Y(n1011) );
  NAND2X1 U1090 ( .A(n124), .B(n1136), .Y(n117) );
  OAI21XL U1091 ( .A0(n152), .A1(n135), .B0(n136), .Y(n134) );
  NOR2X1 U1092 ( .A(n393), .B(n392), .Y(n112) );
  NAND2X1 U1093 ( .A(n453), .B(n461), .Y(n221) );
  OAI21X1 U1094 ( .A0(n156), .A1(n126), .B0(n127), .Y(n125) );
  CLKINVX1 U1095 ( .A(n131), .Y(n129) );
  NOR2X2 U1096 ( .A(n155), .B(n126), .Y(n124) );
  OAI21X1 U1097 ( .A0(n118), .A1(n112), .B0(n113), .Y(n111) );
  OAI21X1 U1098 ( .A0(n346), .A1(n334), .B0(n335), .Y(n333) );
  NAND2X1 U1099 ( .A(n336), .B(n1138), .Y(n334) );
  AOI21X1 U1100 ( .A0(n336), .A1(n342), .B0(n337), .Y(n335) );
  CLKINVX1 U1101 ( .A(n339), .Y(n337) );
  CLKINVX1 U1102 ( .A(n299), .Y(n297) );
  XOR2X2 U1103 ( .A(n1157), .B(n1145), .Y(product[30]) );
  NOR2X1 U1104 ( .A(n557), .B(n565), .Y(n287) );
  NAND2X1 U1105 ( .A(n1164), .B(n1165), .Y(n1167) );
  NAND2X1 U1106 ( .A(n240), .B(n77), .Y(n1166) );
  XOR2X1 U1107 ( .A(n161), .B(n69), .Y(product[29]) );
  CLKXOR2X2 U1108 ( .A(n141), .B(n67), .Y(product[31]) );
  NOR2X1 U1109 ( .A(n497), .B(n508), .Y(n252) );
  NAND2X1 U1110 ( .A(n389), .B(n353), .Y(n96) );
  XNOR2X2 U1111 ( .A(n1189), .B(n82), .Y(product[16]) );
  XNOR2X1 U1112 ( .A(n311), .B(n88), .Y(product[10]) );
  NAND2X2 U1113 ( .A(n1155), .B(n1156), .Y(product[12]) );
  NAND2X1 U1114 ( .A(n1193), .B(n86), .Y(n1155) );
  NAND2X1 U1115 ( .A(n1153), .B(n1154), .Y(n1156) );
  NAND2X1 U1116 ( .A(n1010), .B(n1030), .Y(n1020) );
  XOR2X1 U1117 ( .A(b[2]), .B(b[3]), .Y(n1010) );
  INVXL U1118 ( .A(n220), .Y(n218) );
  OAI22X1 U1119 ( .A0(n916), .A1(n24), .B0(n915), .B1(n22), .Y(n737) );
  XNOR2XL U1120 ( .A(n986), .B(n49), .Y(n824) );
  XNOR2XL U1121 ( .A(n985), .B(n49), .Y(n823) );
  XNOR2X1 U1122 ( .A(n997), .B(n49), .Y(n835) );
  CLKBUFX3 U1123 ( .A(b[18]), .Y(n1133) );
  OAI22X1 U1124 ( .A0(n968), .A1(n6), .B0(n967), .B1(n3), .Y(n789) );
  OAI22XL U1125 ( .A0(n916), .A1(n22), .B0(n917), .B1(n24), .Y(n738) );
  OR2XL U1126 ( .A(n918), .B(n24), .Y(n1175) );
  OAI22XL U1127 ( .A0(n918), .A1(n22), .B0(n919), .B1(n24), .Y(n740) );
  AO21X1 U1128 ( .A0(n24), .A1(n22), .B0(n913), .Y(n734) );
  OAI22XL U1129 ( .A0(n974), .A1(n1031), .B0(n975), .B1(n1021), .Y(n796) );
  INVX3 U1130 ( .A(b[0]), .Y(n1031) );
  NAND2X2 U1131 ( .A(n1004), .B(n1024), .Y(n1014) );
  OR2X1 U1132 ( .A(n413), .B(n409), .Y(n1134) );
  OR2X2 U1133 ( .A(n576), .B(n583), .Y(n1135) );
  OAI21X2 U1134 ( .A0(n167), .A1(n103), .B0(n104), .Y(n102) );
  OR2X1 U1135 ( .A(n395), .B(n394), .Y(n1136) );
  OR2X1 U1136 ( .A(n610), .B(n614), .Y(n1137) );
  CLKBUFX3 U1137 ( .A(b[9]), .Y(n25) );
  OR2X1 U1138 ( .A(n621), .B(n785), .Y(n1138) );
  OR2X1 U1139 ( .A(n400), .B(n396), .Y(n1139) );
  OR2X2 U1140 ( .A(n584), .B(n591), .Y(n1140) );
  INVX1 U1141 ( .A(n156), .Y(n154) );
  OR2X1 U1142 ( .A(n615), .B(n616), .Y(n1141) );
  CLKBUFX3 U1143 ( .A(n1031), .Y(n3) );
  OR2XL U1144 ( .A(n786), .B(n623), .Y(n1142) );
  NAND2X2 U1145 ( .A(n1169), .B(n1134), .Y(n155) );
  OR2X1 U1146 ( .A(n427), .B(n434), .Y(n1143) );
  OR2X1 U1147 ( .A(n391), .B(n634), .Y(n1144) );
  NAND2X1 U1148 ( .A(n1011), .B(n1031), .Y(n1021) );
  XNOR2X2 U1149 ( .A(b[14]), .B(b[13]), .Y(n1024) );
  BUFX4 U1150 ( .A(n1014), .Y(n47) );
  NOR2X1 U1151 ( .A(n605), .B(n609), .Y(n320) );
  BUFX4 U1152 ( .A(n1017), .Y(n30) );
  NOR2X2 U1153 ( .A(n220), .B(n213), .Y(n211) );
  OR2X1 U1154 ( .A(n414), .B(n420), .Y(n1169) );
  NOR2X1 U1155 ( .A(n404), .B(n408), .Y(n146) );
  INVX1 U1156 ( .A(n228), .Y(n226) );
  NOR2X1 U1157 ( .A(n617), .B(n620), .Y(n338) );
  AND2X2 U1158 ( .A(n145), .B(n147), .Y(n1145) );
  NAND2X2 U1159 ( .A(n1003), .B(n1023), .Y(n1013) );
  AND2X2 U1160 ( .A(n357), .B(n113), .Y(n1146) );
  NOR2X1 U1161 ( .A(n453), .B(n461), .Y(n220) );
  NOR2X1 U1162 ( .A(n435), .B(n442), .Y(n202) );
  CLKINVX1 U1163 ( .A(n202), .Y(n200) );
  NOR2X1 U1164 ( .A(n522), .B(n534), .Y(n267) );
  NOR2X1 U1165 ( .A(n426), .B(n421), .Y(n178) );
  CLKINVX1 U1166 ( .A(n178), .Y(n176) );
  CLKINVX1 U1167 ( .A(n1147), .Y(n1148) );
  XNOR2X1 U1168 ( .A(a[1]), .B(n43), .Y(n856) );
  BUFX2 U1169 ( .A(n1019), .Y(n17) );
  ADDFX2 U1170 ( .A(n717), .B(n449), .CI(n671), .CO(n439), .S(n440) );
  NAND2X2 U1171 ( .A(n473), .B(n483), .Y(n239) );
  AOI21X1 U1172 ( .A0(n201), .A1(n187), .B0(n190), .Y(n186) );
  NAND2X2 U1173 ( .A(n1008), .B(n1028), .Y(n1018) );
  XNOR2X2 U1174 ( .A(b[6]), .B(b[5]), .Y(n1028) );
  NAND2X2 U1175 ( .A(n1002), .B(n1022), .Y(n1012) );
  XNOR2X2 U1176 ( .A(n1133), .B(b[17]), .Y(n1022) );
  XNOR2X1 U1177 ( .A(n986), .B(n19), .Y(n914) );
  INVX3 U1178 ( .A(n281), .Y(n1147) );
  OAI21X1 U1179 ( .A0(n174), .A1(n203), .B0(n175), .Y(n173) );
  NAND2X2 U1180 ( .A(n1143), .B(n176), .Y(n174) );
  CMPR42X2 U1181 ( .A(n466), .B(n659), .C(n673), .D(n703), .ICI(n463), .S(n456), .ICO(n454), .CO(n455) );
  AOI21X4 U1182 ( .A0(n190), .A1(n176), .B0(n177), .Y(n175) );
  NAND2X4 U1183 ( .A(n1132), .B(n229), .Y(n227) );
  NOR2X2 U1184 ( .A(n238), .B(n231), .Y(n229) );
  XNOR2X2 U1185 ( .A(n986), .B(n25), .Y(n896) );
  OAI21X1 U1186 ( .A0(n205), .A1(n254), .B0(n206), .Y(n204) );
  NAND2XL U1187 ( .A(n225), .B(n211), .Y(n205) );
  CMPR42X2 U1188 ( .A(n514), .B(n503), .C(n511), .D(n500), .ICI(n507), .S(n497), .ICO(n495), .CO(n496) );
  OAI22X1 U1189 ( .A0(n979), .A1(n3), .B0(n980), .B1(n6), .Y(n801) );
  XNOR2X1 U1190 ( .A(a[3]), .B(n1), .Y(n980) );
  XNOR2X1 U1191 ( .A(n993), .B(n31), .Y(n885) );
  XNOR2X1 U1192 ( .A(n985), .B(n7), .Y(n949) );
  OAI21X1 U1193 ( .A0(n309), .A1(n313), .B0(n310), .Y(n308) );
  XNOR2X1 U1194 ( .A(a[3]), .B(n37), .Y(n872) );
  CLKBUFX8 U1195 ( .A(b[13]), .Y(n37) );
  OAI21X2 U1196 ( .A0(n194), .A1(n254), .B0(n195), .Y(n193) );
  NAND2XL U1197 ( .A(n225), .B(n196), .Y(n194) );
  AOI21X4 U1198 ( .A0(n248), .A1(n229), .B0(n230), .Y(n228) );
  OAI21X1 U1199 ( .A0(n231), .A1(n239), .B0(n232), .Y(n230) );
  OAI21X1 U1200 ( .A0(n292), .A1(n290), .B0(n291), .Y(n289) );
  INVX1 U1201 ( .A(n293), .Y(n292) );
  CMPR42X2 U1202 ( .A(n532), .B(n542), .C(n772), .D(n664), .ICI(n756), .S(n528), .ICO(n526), .CO(n527) );
  XNOR2X1 U1203 ( .A(n987), .B(n19), .Y(n915) );
  XNOR2X1 U1204 ( .A(n987), .B(n31), .Y(n879) );
  CMPR42X2 U1205 ( .A(n1125), .B(n1126), .C(n738), .D(n506), .ICI(n510), .S(
        n500), .ICO(n498), .CO(n499) );
  XNOR2X1 U1206 ( .A(n987), .B(n37), .Y(n861) );
  XNOR2X1 U1207 ( .A(n993), .B(n25), .Y(n903) );
  XNOR2X1 U1208 ( .A(n987), .B(n25), .Y(n897) );
  OAI22X1 U1209 ( .A0(n866), .A1(n40), .B0(n867), .B1(n41), .Y(n690) );
  OAI22X1 U1210 ( .A0(n868), .A1(n41), .B0(n867), .B1(n39), .Y(n691) );
  OAI22X1 U1211 ( .A0(n861), .A1(n41), .B0(n860), .B1(n40), .Y(n684) );
  OAI22X1 U1212 ( .A0(n862), .A1(n41), .B0(n861), .B1(n40), .Y(n685) );
  XNOR2X1 U1213 ( .A(n988), .B(n13), .Y(n934) );
  OAI21X1 U1214 ( .A0(n314), .A1(n312), .B0(n313), .Y(n311) );
  ADDFHX2 U1215 ( .A(n494), .B(n753), .CI(n721), .CO(n491), .S(n492) );
  OAI22X4 U1216 ( .A0(n846), .A1(n47), .B0(n845), .B1(n46), .Y(n670) );
  OAI21X1 U1217 ( .A0(n216), .A1(n254), .B0(n217), .Y(n215) );
  INVX8 U1218 ( .A(n255), .Y(n254) );
  AOI21XL U1219 ( .A0(n226), .A1(n218), .B0(n219), .Y(n217) );
  XOR2X4 U1220 ( .A(n123), .B(n65), .Y(product[33]) );
  XNOR2X1 U1221 ( .A(a[1]), .B(n49), .Y(n838) );
  OAI22X1 U1222 ( .A0(n942), .A1(n15), .B0(n943), .B1(n17), .Y(n764) );
  XNOR2X1 U1223 ( .A(n988), .B(n19), .Y(n916) );
  CLKINVX3 U1224 ( .A(n306), .Y(n305) );
  AOI21X2 U1225 ( .A0(n307), .A1(n315), .B0(n308), .Y(n306) );
  XNOR2X4 U1226 ( .A(n289), .B(n84), .Y(product[14]) );
  OAI22X1 U1227 ( .A0(n933), .A1(n18), .B0(n932), .B1(n16), .Y(n754) );
  XOR2X4 U1228 ( .A(n109), .B(n63), .Y(product[35]) );
  XNOR2X2 U1229 ( .A(a[3]), .B(n25), .Y(n908) );
  XNOR2X1 U1230 ( .A(a[1]), .B(n37), .Y(n874) );
  XNOR2X4 U1231 ( .A(n215), .B(n74), .Y(product[24]) );
  OAI22X2 U1232 ( .A0(n835), .A1(n52), .B0(n836), .B1(n1013), .Y(n493) );
  XNOR2X1 U1233 ( .A(a[3]), .B(n49), .Y(n836) );
  CLKBUFX3 U1234 ( .A(a[8]), .Y(n993) );
  BUFX12 U1235 ( .A(a[16]), .Y(n985) );
  AOI21X1 U1236 ( .A0(n283), .A1(n263), .B0(n264), .Y(n262) );
  XNOR2X1 U1237 ( .A(n995), .B(n49), .Y(n833) );
  OR2X4 U1238 ( .A(n984), .B(n3), .Y(n1149) );
  OR2X1 U1239 ( .A(n6), .B(n1041), .Y(n1150) );
  NAND2X6 U1240 ( .A(n1149), .B(n1150), .Y(n633) );
  NAND2BXL U1241 ( .AN(n61), .B(n1), .Y(n984) );
  INVXL U1242 ( .A(n1), .Y(n1041) );
  NOR2X2 U1243 ( .A(n804), .B(n633), .Y(n354) );
  NAND2X6 U1244 ( .A(n804), .B(n633), .Y(n355) );
  XOR2X4 U1245 ( .A(n132), .B(n66), .Y(product[32]) );
  XNOR2X1 U1246 ( .A(n989), .B(n43), .Y(n845) );
  BUFX12 U1247 ( .A(a[12]), .Y(n989) );
  XNOR2X4 U1248 ( .A(n204), .B(n73), .Y(product[25]) );
  OR2XL U1249 ( .A(n836), .B(n52), .Y(n1151) );
  OR2X1 U1250 ( .A(n837), .B(n1013), .Y(n1152) );
  NAND2X1 U1251 ( .A(n1151), .B(n1152), .Y(n662) );
  CMPR42X2 U1252 ( .A(n662), .B(n770), .C(n677), .D(n722), .ICI(n518), .S(n506), .ICO(n504), .CO(n505) );
  INVX3 U1253 ( .A(n1193), .Y(n1153) );
  CLKINVX1 U1254 ( .A(n86), .Y(n1154) );
  AO21X1 U1255 ( .A0(n305), .A1(n1140), .B0(n302), .Y(n1193) );
  AO21XL U1256 ( .A0(n1177), .A1(n153), .B0(n154), .Y(n1157) );
  NAND2XL U1257 ( .A(n994), .B(n49), .Y(n1160) );
  NAND2X1 U1258 ( .A(n1158), .B(n1159), .Y(n1161) );
  NAND2X1 U1259 ( .A(n1160), .B(n1161), .Y(n832) );
  INVXL U1260 ( .A(n994), .Y(n1158) );
  INVXL U1261 ( .A(n49), .Y(n1159) );
  BUFX12 U1262 ( .A(a[7]), .Y(n994) );
  OAI22X1 U1263 ( .A0(n832), .A1(n1013), .B0(n831), .B1(n52), .Y(n658) );
  OAI22X1 U1264 ( .A0(n833), .A1(n1013), .B0(n832), .B1(n52), .Y(n659) );
  AOI2BB1X4 U1265 ( .A0N(n181), .A1N(n254), .B0(n1163), .Y(n1162) );
  CLKINVX20 U1266 ( .A(n1162), .Y(n180) );
  AO21XL U1267 ( .A0(n226), .A1(n183), .B0(n184), .Y(n1163) );
  XNOR2X4 U1268 ( .A(n180), .B(n71), .Y(product[27]) );
  XNOR2X1 U1269 ( .A(n995), .B(n55), .Y(n815) );
  BUFX12 U1270 ( .A(a[6]), .Y(n995) );
  CLKINVX4 U1271 ( .A(n240), .Y(n1164) );
  CLKINVX1 U1272 ( .A(n77), .Y(n1165) );
  OAI21X4 U1273 ( .A0(n254), .A1(n241), .B0(n246), .Y(n240) );
  NAND2XL U1274 ( .A(n236), .B(n239), .Y(n77) );
  ADDHX2 U1275 ( .A(n748), .B(n764), .CO(n601), .S(n602) );
  XOR2X4 U1276 ( .A(n1168), .B(n78), .Y(product[20]) );
  OA21XL U1277 ( .A0(n254), .A1(n252), .B0(n253), .Y(n1168) );
  CLKINVX2 U1278 ( .A(n227), .Y(n225) );
  NOR2X2 U1279 ( .A(n174), .B(n202), .Y(n172) );
  NAND2X4 U1280 ( .A(n1170), .B(n1171), .Y(n753) );
  OR2XL U1281 ( .A(n931), .B(n16), .Y(n1171) );
  OR2X1 U1282 ( .A(n932), .B(n18), .Y(n1170) );
  NAND2XL U1283 ( .A(n992), .B(n25), .Y(n1173) );
  CMPR42X2 U1284 ( .A(n640), .B(n668), .C(n416), .D(n423), .ICI(n419), .S(n414), .ICO(n412), .CO(n413) );
  CMPR42X2 U1285 ( .A(n1124), .B(n669), .C(n429), .D(n424), .ICI(n425), .S(
        n421), .ICO(n419), .CO(n420) );
  XNOR2X1 U1286 ( .A(n986), .B(n37), .Y(n860) );
  NAND2X1 U1287 ( .A(n225), .B(n183), .Y(n181) );
  NAND2X1 U1288 ( .A(n225), .B(n218), .Y(n216) );
  NAND2X1 U1289 ( .A(n1172), .B(n1037), .Y(n1174) );
  CLKBUFX2 U1290 ( .A(n1029), .Y(n16) );
  CLKBUFX2 U1291 ( .A(n1019), .Y(n18) );
  XNOR2X1 U1292 ( .A(n985), .B(n13), .Y(n931) );
  INVX1 U1293 ( .A(n1177), .Y(n167) );
  NAND2X1 U1294 ( .A(n592), .B(n597), .Y(n310) );
  NOR2X2 U1295 ( .A(n803), .B(n787), .Y(n352) );
  BUFX8 U1296 ( .A(a[10]), .Y(n991) );
  INVXL U1297 ( .A(n992), .Y(n1172) );
  AO21XL U1298 ( .A0(n1177), .A1(n115), .B0(n116), .Y(n1181) );
  ADDHX1 U1299 ( .A(n766), .B(n782), .CO(n611), .S(n612) );
  OR2XL U1300 ( .A(n917), .B(n22), .Y(n1176) );
  ADDFHX1 U1301 ( .A(n649), .B(n531), .CI(n739), .CO(n516), .S(n517) );
  XNOR2X1 U1302 ( .A(n989), .B(n25), .Y(n899) );
  BUFX12 U1303 ( .A(a[9]), .Y(n992) );
  AOI21X1 U1304 ( .A0(n111), .A1(n1144), .B0(n106), .Y(n104) );
  OAI22X1 U1305 ( .A0(n884), .A1(n36), .B0(n883), .B1(n34), .Y(n706) );
  OR2X4 U1306 ( .A(n982), .B(n3), .Y(n1179) );
  OR2X4 U1307 ( .A(n983), .B(n6), .Y(n1180) );
  NAND2X1 U1308 ( .A(n1182), .B(n1183), .Y(n1185) );
  CLKBUFX2 U1309 ( .A(n1028), .Y(n22) );
  CLKBUFX2 U1310 ( .A(n1018), .Y(n24) );
  OAI2BB1X4 U1311 ( .A0N(n168), .A1N(n255), .B0(n1178), .Y(n1177) );
  OA21XL U1312 ( .A0(n228), .A1(n170), .B0(n171), .Y(n1178) );
  NAND2X1 U1313 ( .A(n110), .B(n1144), .Y(n103) );
  OAI22X1 U1314 ( .A0(n890), .A1(n34), .B0(n891), .B1(n35), .Y(n713) );
  NAND2BXL U1315 ( .AN(n354), .B(n355), .Y(n97) );
  OAI22XL U1316 ( .A0(n964), .A1(n11), .B0(n963), .B1(n9), .Y(n785) );
  NAND2X1 U1317 ( .A(n615), .B(n616), .Y(n332) );
  XNOR2X1 U1318 ( .A(n986), .B(n7), .Y(n950) );
  XNOR2X1 U1319 ( .A(n994), .B(n37), .Y(n868) );
  ADDFX2 U1320 ( .A(n602), .B(n629), .CI(n606), .CO(n599), .S(n600) );
  NAND2XL U1321 ( .A(a[3]), .B(n43), .Y(n1184) );
  NAND2X2 U1322 ( .A(n1184), .B(n1185), .Y(n854) );
  INVXL U1323 ( .A(a[3]), .Y(n1182) );
  NAND2X4 U1324 ( .A(n1179), .B(n1180), .Y(n804) );
  XNOR2XL U1325 ( .A(n61), .B(n1), .Y(n983) );
  NOR2X2 U1326 ( .A(n209), .B(n198), .Y(n196) );
  AOI21XL U1327 ( .A0(n226), .A1(n211), .B0(n212), .Y(n206) );
  CLKINVX8 U1328 ( .A(n102), .Y(n101) );
  NAND2X1 U1329 ( .A(n462), .B(n472), .Y(n232) );
  NOR2X2 U1330 ( .A(n509), .B(n521), .Y(n260) );
  AOI21X2 U1331 ( .A0(n333), .A1(n1141), .B0(n330), .Y(n328) );
  NAND2XL U1332 ( .A(n1140), .B(n304), .Y(n87) );
  CMPR42X1 U1333 ( .A(n680), .B(n550), .C(n710), .D(n741), .ICI(n551), .S(n538), .ICO(n536), .CO(n537) );
  OR2X4 U1334 ( .A(n855), .B(n47), .Y(n1187) );
  NAND2X2 U1335 ( .A(n1186), .B(n1187), .Y(n679) );
  OR2X4 U1336 ( .A(n854), .B(n1024), .Y(n1186) );
  CMPR32X2 U1337 ( .A(n450), .B(n687), .C(n457), .CO(n447), .S(n448) );
  XNOR2XL U1338 ( .A(n993), .B(n37), .Y(n867) );
  XOR2X1 U1339 ( .A(b[16]), .B(b[17]), .Y(n1003) );
  CLKBUFX3 U1340 ( .A(b[1]), .Y(n1) );
  CLKXOR2X1 U1341 ( .A(b[10]), .B(b[11]), .Y(n1006) );
  CLKXOR2X1 U1342 ( .A(b[6]), .B(b[7]), .Y(n1008) );
  CLKBUFX4 U1343 ( .A(b[19]), .Y(n55) );
  CLKBUFX3 U1344 ( .A(b[15]), .Y(n43) );
  XOR2X4 U1345 ( .A(n1181), .B(n1146), .Y(product[34]) );
  INVX1 U1346 ( .A(n43), .Y(n1183) );
  NAND2X1 U1347 ( .A(n1132), .B(n236), .Y(n234) );
  OAI21X2 U1348 ( .A0(n249), .A1(n253), .B0(n250), .Y(n248) );
  AOI21X1 U1349 ( .A0(n244), .A1(n236), .B0(n237), .Y(n235) );
  NAND2X1 U1350 ( .A(n200), .B(n187), .Y(n185) );
  BUFX20 U1351 ( .A(n101), .Y(\product[39] ) );
  INVXL U1352 ( .A(n252), .Y(n372) );
  INVX3 U1353 ( .A(n320), .Y(n318) );
  OA21X4 U1354 ( .A0(n287), .A1(n291), .B0(n288), .Y(n1192) );
  NAND2X1 U1355 ( .A(n376), .B(n282), .Y(n83) );
  INVXL U1356 ( .A(n1148), .Y(n376) );
  OAI21X2 U1357 ( .A0(n276), .A1(n282), .B0(n277), .Y(n275) );
  INVXL U1358 ( .A(n312), .Y(n382) );
  NAND2X2 U1359 ( .A(n605), .B(n609), .Y(n321) );
  NAND2X1 U1360 ( .A(n1135), .B(n1140), .Y(n294) );
  NAND2X1 U1361 ( .A(n566), .B(n575), .Y(n291) );
  NAND2X1 U1362 ( .A(n610), .B(n614), .Y(n326) );
  INVX3 U1363 ( .A(n304), .Y(n302) );
  OR2X4 U1364 ( .A(n961), .B(n11), .Y(n1196) );
  NAND2X2 U1365 ( .A(n1195), .B(n1196), .Y(n782) );
  OAI22XL U1366 ( .A0(n959), .A1(n11), .B0(n958), .B1(n9), .Y(n780) );
  OAI22XL U1367 ( .A0(n887), .A1(n34), .B0(n888), .B1(n35), .Y(n710) );
  OAI22X1 U1368 ( .A0(n814), .A1(n59), .B0(n813), .B1(n57), .Y(n642) );
  CMPR42X1 U1369 ( .A(n793), .B(n761), .C(n581), .D(n714), .ICI(n777), .S(n579), .ICO(n577), .CO(n578) );
  OAI22XL U1370 ( .A0(n1123), .A1(n12), .B0(n955), .B1(n9), .Y(n777) );
  OAI22X2 U1371 ( .A0(n878), .A1(n36), .B0(n877), .B1(n34), .Y(n431) );
  XNOR2XL U1372 ( .A(n788), .B(n679), .Y(n532) );
  BUFX8 U1373 ( .A(a[14]), .Y(n987) );
  XNOR2X1 U1374 ( .A(n992), .B(n31), .Y(n884) );
  XNOR2X1 U1375 ( .A(n992), .B(n37), .Y(n866) );
  NAND2BXL U1376 ( .AN(n61), .B(n25), .Y(n912) );
  XNOR2X1 U1377 ( .A(n994), .B(n31), .Y(n886) );
  XNOR2X1 U1378 ( .A(n987), .B(n13), .Y(n933) );
  XNOR2X1 U1379 ( .A(n991), .B(n43), .Y(n847) );
  BUFX8 U1380 ( .A(a[4]), .Y(n997) );
  CLKBUFX4 U1381 ( .A(b[5]), .Y(n13) );
  XNOR2X1 U1382 ( .A(b[2]), .B(b[1]), .Y(n1030) );
  XNOR2X1 U1383 ( .A(b[8]), .B(b[7]), .Y(n1027) );
  CLKBUFX4 U1384 ( .A(b[7]), .Y(n19) );
  INVX1 U1385 ( .A(n1132), .Y(n241) );
  NOR2XL U1386 ( .A(n272), .B(n265), .Y(n263) );
  INVXL U1387 ( .A(n273), .Y(n271) );
  XOR2X4 U1388 ( .A(n1188), .B(n75), .Y(product[23]) );
  OA21XL U1389 ( .A0(n254), .A1(n227), .B0(n228), .Y(n1188) );
  OAI21X4 U1390 ( .A0(n284), .A1(n256), .B0(n257), .Y(n255) );
  NAND2XL U1391 ( .A(n372), .B(n253), .Y(n79) );
  AO21XL U1392 ( .A0(n283), .A1(n376), .B0(n280), .Y(n1189) );
  NAND2XL U1393 ( .A(n373), .B(n261), .Y(n80) );
  INVXL U1394 ( .A(n239), .Y(n237) );
  CLKINVX1 U1395 ( .A(n211), .Y(n209) );
  NOR2XL U1396 ( .A(n155), .B(n144), .Y(n142) );
  OAI21X2 U1397 ( .A0(n316), .A1(n328), .B0(n317), .Y(n315) );
  AOI21X2 U1398 ( .A0(n318), .A1(n324), .B0(n319), .Y(n317) );
  NAND2X2 U1399 ( .A(n318), .B(n1137), .Y(n316) );
  OA21X4 U1400 ( .A0(n1190), .A1(n1191), .B0(n1192), .Y(n284) );
  OR2X2 U1401 ( .A(n287), .B(n290), .Y(n1191) );
  NOR2X2 U1402 ( .A(n1148), .B(n276), .Y(n274) );
  AOI21XL U1403 ( .A0(n327), .A1(n1137), .B0(n324), .Y(n322) );
  NAND2XL U1404 ( .A(n382), .B(n313), .Y(n89) );
  NAND2XL U1405 ( .A(n377), .B(n288), .Y(n84) );
  INVXL U1406 ( .A(n287), .Y(n377) );
  NAND2XL U1407 ( .A(n1138), .B(n344), .Y(n94) );
  INVXL U1408 ( .A(n309), .Y(n381) );
  OAI21X4 U1409 ( .A0(n139), .A1(n147), .B0(n140), .Y(n138) );
  OAI21X2 U1410 ( .A0(n213), .A1(n221), .B0(n214), .Y(n212) );
  AOI21X2 U1411 ( .A0(n125), .A1(n1136), .B0(n120), .Y(n118) );
  AOI21X2 U1412 ( .A0(n163), .A1(n1134), .B0(n158), .Y(n156) );
  NOR2X4 U1413 ( .A(n146), .B(n139), .Y(n137) );
  INVXL U1414 ( .A(n203), .Y(n201) );
  INVXL U1415 ( .A(n282), .Y(n280) );
  OAI21X4 U1416 ( .A0(n306), .A1(n294), .B0(n295), .Y(n293) );
  CMPR42X2 U1417 ( .A(n527), .B(n515), .C(n524), .D(n512), .ICI(n520), .S(n509), .ICO(n507), .CO(n508) );
  CMPR42X2 U1418 ( .A(n558), .B(n552), .C(n559), .D(n549), .ICI(n555), .S(n546), .ICO(n544), .CO(n545) );
  CMPR42X2 U1419 ( .A(n536), .B(n528), .C(n537), .D(n525), .ICI(n533), .S(n522), .ICO(n520), .CO(n521) );
  NOR2X1 U1420 ( .A(n546), .B(n556), .Y(n281) );
  NOR2X1 U1421 ( .A(n598), .B(n604), .Y(n312) );
  INVXL U1422 ( .A(n352), .Y(n389) );
  AO21XL U1423 ( .A0(n345), .A1(n1138), .B0(n342), .Y(n1194) );
  ADDHX1 U1424 ( .A(n730), .B(n746), .CO(n588), .S(n589) );
  OAI22X2 U1425 ( .A0(n924), .A1(n21), .B0(n925), .B1(n23), .Y(n746) );
  ADDHX1 U1426 ( .A(n696), .B(n711), .CO(n553), .S(n554) );
  OAI22X1 U1427 ( .A0(n872), .A1(n39), .B0(n873), .B1(n41), .Y(n696) );
  OAI22X1 U1428 ( .A0(n962), .A1(n9), .B0(n963), .B1(n11), .Y(n784) );
  ADDHX1 U1429 ( .A(n713), .B(n728), .CO(n572), .S(n573) );
  CMPR32X2 U1430 ( .A(n694), .B(n740), .C(n625), .CO(n529), .S(n530) );
  CMPR42X2 U1431 ( .A(n759), .B(n567), .C(n568), .D(n560), .ICI(n564), .S(n557), .ICO(n555), .CO(n556) );
  CMPR42X2 U1432 ( .A(n732), .B(n780), .C(n796), .D(n600), .ICI(n603), .S(n598), .ICO(n596), .CO(n597) );
  CMPR32X2 U1433 ( .A(n801), .B(n769), .C(n622), .CO(n620), .S(n621) );
  NOR2BXL U1434 ( .AN(n61), .B(n15), .Y(n769) );
  OAI22X1 U1435 ( .A0(n816), .A1(n57), .B0(n817), .B1(n59), .Y(n645) );
  ADDFX2 U1436 ( .A(n695), .B(n789), .CI(n665), .CO(n542), .S(n543) );
  NOR2BXL U1437 ( .AN(n61), .B(n52), .Y(n665) );
  AO21XL U1438 ( .A0(n41), .A1(n40), .B0(n859), .Y(n683) );
  AO21XL U1439 ( .A0(n30), .A1(n28), .B0(n895), .Y(n717) );
  ADDFX1 U1440 ( .A(n646), .B(n493), .CI(n752), .CO(n480), .S(n481) );
  AO21XL U1441 ( .A0(n18), .A1(n16), .B0(n931), .Y(n752) );
  INVXL U1442 ( .A(n449), .Y(n450) );
  INVXL U1443 ( .A(n493), .Y(n494) );
  NOR2BXL U1444 ( .AN(n61), .B(n1024), .Y(n682) );
  CMPR42X2 U1445 ( .A(n504), .B(n691), .C(n647), .D(n492), .ICI(n505), .S(n490), .ICO(n488), .CO(n489) );
  CMPR42X2 U1446 ( .A(n660), .B(n477), .C(n1128), .D(n719), .ICI(n478), .S(
        n465), .ICO(n463), .CO(n464) );
  CMPR42X2 U1447 ( .A(n643), .B(n686), .C(n445), .D(n438), .ICI(n441), .S(n435), .ICO(n433), .CO(n434) );
  OAI22X1 U1448 ( .A0(n817), .A1(n57), .B0(n818), .B1(n59), .Y(n469) );
  ADDFXL U1449 ( .A(n650), .B(n397), .CI(n635), .CO(n393), .S(n394) );
  AO21XL U1450 ( .A0(n54), .A1(n52), .B0(n823), .Y(n650) );
  OAI22XL U1451 ( .A0(n824), .A1(n54), .B0(n823), .B1(n52), .Y(n397) );
  OAI22X1 U1452 ( .A0(n806), .A1(n60), .B0(n805), .B1(n58), .Y(n391) );
  AO21XL U1453 ( .A0(n60), .A1(n58), .B0(n805), .Y(n634) );
  XNOR2XL U1454 ( .A(n992), .B(n7), .Y(n956) );
  ADDFX2 U1455 ( .A(n573), .B(n776), .CI(n627), .CO(n570), .S(n571) );
  NAND2BXL U1456 ( .AN(n61), .B(n7), .Y(n966) );
  NAND2BXL U1457 ( .AN(n61), .B(n13), .Y(n948) );
  NAND2BXL U1458 ( .AN(n61), .B(n49), .Y(n840) );
  NAND2BXL U1459 ( .AN(n61), .B(n19), .Y(n930) );
  NAND2BXL U1460 ( .AN(n61), .B(n37), .Y(n876) );
  OAI22X2 U1461 ( .A0(n966), .A1(n9), .B0(n12), .B1(n1040), .Y(n632) );
  OAI22X2 U1462 ( .A0(n948), .A1(n16), .B0(n18), .B1(n1039), .Y(n631) );
  XNOR2XL U1463 ( .A(n991), .B(n13), .Y(n937) );
  XNOR2XL U1464 ( .A(n989), .B(n1), .Y(n971) );
  XNOR2XL U1465 ( .A(n989), .B(n7), .Y(n953) );
  XNOR2XL U1466 ( .A(n994), .B(n55), .Y(n814) );
  XNOR2XL U1467 ( .A(n994), .B(n13), .Y(n940) );
  XNOR2XL U1468 ( .A(n994), .B(n25), .Y(n904) );
  XNOR2XL U1469 ( .A(n994), .B(n19), .Y(n922) );
  XNOR2XL U1470 ( .A(a[3]), .B(n31), .Y(n890) );
  XNOR2XL U1471 ( .A(a[3]), .B(n7), .Y(n962) );
  XNOR2XL U1472 ( .A(n994), .B(n43), .Y(n850) );
  XNOR2XL U1473 ( .A(n992), .B(n13), .Y(n938) );
  XNOR2XL U1474 ( .A(n992), .B(n55), .Y(n812) );
  XNOR2XL U1475 ( .A(a[1]), .B(n31), .Y(n892) );
  XNOR2XL U1476 ( .A(n992), .B(n43), .Y(n848) );
  XNOR2XL U1477 ( .A(n985), .B(n19), .Y(n913) );
  XNOR2XL U1478 ( .A(n61), .B(n25), .Y(n911) );
  XNOR2XL U1479 ( .A(n61), .B(n19), .Y(n929) );
  XNOR2XL U1480 ( .A(n61), .B(n43), .Y(n857) );
  XNOR2XL U1481 ( .A(n61), .B(n49), .Y(n839) );
  XNOR2XL U1482 ( .A(n61), .B(n55), .Y(n821) );
  NAND2BXL U1483 ( .AN(n61), .B(n31), .Y(n894) );
  NAND2BXL U1484 ( .AN(n61), .B(n43), .Y(n858) );
  NAND2BXL U1485 ( .AN(n61), .B(n55), .Y(n822) );
  XNOR2XL U1486 ( .A(n991), .B(n55), .Y(n811) );
  XNOR2XL U1487 ( .A(n989), .B(n49), .Y(n827) );
  XNOR2XL U1488 ( .A(n993), .B(n55), .Y(n813) );
  XNOR2XL U1489 ( .A(n989), .B(n31), .Y(n881) );
  XNOR2XL U1490 ( .A(n989), .B(n55), .Y(n809) );
  XNOR2XL U1491 ( .A(n993), .B(n19), .Y(n921) );
  XNOR2XL U1492 ( .A(n991), .B(n37), .Y(n865) );
  XNOR2XL U1493 ( .A(n991), .B(n49), .Y(n829) );
  XNOR2XL U1494 ( .A(n993), .B(n49), .Y(n831) );
  XNOR2XL U1495 ( .A(n993), .B(n43), .Y(n849) );
  XNOR2XL U1496 ( .A(n987), .B(n55), .Y(n807) );
  XNOR2XL U1497 ( .A(n987), .B(n43), .Y(n843) );
  XNOR2XL U1498 ( .A(n987), .B(n49), .Y(n825) );
  XNOR2XL U1499 ( .A(n988), .B(n55), .Y(n808) );
  XNOR2XL U1500 ( .A(n988), .B(n37), .Y(n862) );
  XNOR2XL U1501 ( .A(n988), .B(n49), .Y(n826) );
  XNOR2XL U1502 ( .A(n990), .B(n55), .Y(n810) );
  XNOR2XL U1503 ( .A(n990), .B(n49), .Y(n828) );
  XNOR2XL U1504 ( .A(n985), .B(n43), .Y(n841) );
  CLKBUFX3 U1505 ( .A(n1030), .Y(n9) );
  CLKBUFX3 U1506 ( .A(n1020), .Y(n11) );
  XNOR2X1 U1507 ( .A(b[10]), .B(b[9]), .Y(n1026) );
  NAND2X4 U1508 ( .A(n1009), .B(n1029), .Y(n1019) );
  NAND2X4 U1509 ( .A(n1006), .B(n1026), .Y(n1016) );
  XNOR2X1 U1510 ( .A(b[12]), .B(b[11]), .Y(n1025) );
  XOR2X4 U1511 ( .A(n1197), .B(n76), .Y(product[22]) );
  OA21XL U1512 ( .A0(n254), .A1(n234), .B0(n235), .Y(n1197) );
  NOR2X1 U1513 ( .A(n209), .B(n185), .Y(n183) );
  CLKINVX1 U1514 ( .A(n246), .Y(n244) );
  CLKINVX1 U1515 ( .A(n248), .Y(n246) );
  CLKINVX1 U1516 ( .A(n155), .Y(n153) );
  NOR2X1 U1517 ( .A(n155), .B(n135), .Y(n133) );
  CLKINVX1 U1518 ( .A(n117), .Y(n115) );
  NOR2X1 U1519 ( .A(n227), .B(n170), .Y(n168) );
  NAND2X1 U1520 ( .A(n211), .B(n172), .Y(n170) );
  NAND2X1 U1521 ( .A(n218), .B(n221), .Y(n75) );
  NAND2X1 U1522 ( .A(n369), .B(n232), .Y(n76) );
  CLKINVX1 U1523 ( .A(n231), .Y(n369) );
  NAND2X1 U1524 ( .A(n258), .B(n274), .Y(n256) );
  NOR2X1 U1525 ( .A(n260), .B(n267), .Y(n258) );
  OAI21XL U1526 ( .A0(n273), .A1(n265), .B0(n268), .Y(n264) );
  CLKINVX1 U1527 ( .A(n221), .Y(n219) );
  OAI21XL U1528 ( .A0(n210), .A1(n185), .B0(n186), .Y(n184) );
  AOI21X1 U1529 ( .A0(n226), .A1(n196), .B0(n197), .Y(n195) );
  OAI21XL U1530 ( .A0(n210), .A1(n198), .B0(n203), .Y(n197) );
  CLKINVX1 U1531 ( .A(n260), .Y(n373) );
  NAND2X1 U1532 ( .A(n266), .B(n268), .Y(n81) );
  AOI21X1 U1533 ( .A0(n283), .A1(n274), .B0(n271), .Y(n269) );
  NAND2X1 U1534 ( .A(n375), .B(n277), .Y(n82) );
  CLKINVX1 U1535 ( .A(n276), .Y(n375) );
  XOR2X1 U1536 ( .A(n254), .B(n79), .Y(product[19]) );
  NAND2X1 U1537 ( .A(n371), .B(n250), .Y(n78) );
  CLKINVX1 U1538 ( .A(n249), .Y(n371) );
  CLKINVX1 U1539 ( .A(n284), .Y(n283) );
  CLKINVX1 U1540 ( .A(n212), .Y(n210) );
  NAND2X1 U1541 ( .A(n137), .B(n1139), .Y(n126) );
  CLKINVX1 U1542 ( .A(n274), .Y(n272) );
  CLKINVX1 U1543 ( .A(n238), .Y(n236) );
  CLKINVX1 U1544 ( .A(n275), .Y(n273) );
  CLKINVX1 U1545 ( .A(n315), .Y(n314) );
  CLKINVX1 U1546 ( .A(n200), .Y(n198) );
  CLKINVX1 U1547 ( .A(n266), .Y(n265) );
  CLKINVX1 U1548 ( .A(n267), .Y(n266) );
  CLKINVX1 U1549 ( .A(n188), .Y(n187) );
  CLKINVX1 U1550 ( .A(n1143), .Y(n188) );
  CLKINVX1 U1551 ( .A(n118), .Y(n116) );
  CLKINVX1 U1552 ( .A(n138), .Y(n136) );
  CLKINVX1 U1553 ( .A(n154), .Y(n152) );
  CLKINVX1 U1554 ( .A(n137), .Y(n135) );
  NOR2X2 U1555 ( .A(n462), .B(n472), .Y(n231) );
  NOR2X2 U1556 ( .A(n484), .B(n496), .Y(n249) );
  AOI21X1 U1557 ( .A0(n172), .A1(n212), .B0(n173), .Y(n171) );
  CLKINVX1 U1558 ( .A(n179), .Y(n177) );
  NAND2X1 U1559 ( .A(n497), .B(n508), .Y(n253) );
  NAND2X1 U1560 ( .A(n484), .B(n496), .Y(n250) );
  XNOR2X1 U1561 ( .A(n1177), .B(n70), .Y(product[28]) );
  NAND2X1 U1562 ( .A(n1169), .B(n165), .Y(n70) );
  NAND2X1 U1563 ( .A(n176), .B(n179), .Y(n71) );
  NAND2X1 U1564 ( .A(n187), .B(n192), .Y(n72) );
  NAND2X1 U1565 ( .A(n200), .B(n203), .Y(n73) );
  NAND2X1 U1566 ( .A(n367), .B(n214), .Y(n74) );
  CLKINVX1 U1567 ( .A(n213), .Y(n367) );
  XNOR2X1 U1568 ( .A(n283), .B(n83), .Y(product[15]) );
  NAND2X1 U1569 ( .A(n381), .B(n310), .Y(n88) );
  XNOR2X1 U1570 ( .A(n327), .B(n91), .Y(product[7]) );
  NAND2X1 U1571 ( .A(n1137), .B(n326), .Y(n91) );
  XNOR2X1 U1572 ( .A(n345), .B(n94), .Y(product[4]) );
  NOR2X1 U1573 ( .A(n309), .B(n312), .Y(n307) );
  CLKINVX1 U1574 ( .A(n321), .Y(n319) );
  NOR2X2 U1575 ( .A(n535), .B(n545), .Y(n276) );
  AOI21X1 U1576 ( .A0(n138), .A1(n1139), .B0(n129), .Y(n127) );
  NAND2X1 U1577 ( .A(n1144), .B(n108), .Y(n63) );
  AOI21X1 U1578 ( .A0(n1177), .A1(n110), .B0(n111), .Y(n109) );
  XOR2X1 U1579 ( .A(n292), .B(n85), .Y(product[13]) );
  NAND2X1 U1580 ( .A(n378), .B(n291), .Y(n85) );
  CLKINVX1 U1581 ( .A(n290), .Y(n378) );
  NAND2X1 U1582 ( .A(n318), .B(n321), .Y(n90) );
  CLKINVX1 U1583 ( .A(n112), .Y(n357) );
  NAND2X1 U1584 ( .A(n1136), .B(n122), .Y(n65) );
  AOI21X1 U1585 ( .A0(n1177), .A1(n124), .B0(n125), .Y(n123) );
  NAND2X1 U1586 ( .A(n360), .B(n140), .Y(n67) );
  AOI21X1 U1587 ( .A0(n1177), .A1(n142), .B0(n143), .Y(n141) );
  CLKINVX1 U1588 ( .A(n139), .Y(n360) );
  NAND2X1 U1589 ( .A(n1134), .B(n160), .Y(n69) );
  AOI21X1 U1590 ( .A0(n1177), .A1(n1169), .B0(n163), .Y(n161) );
  NAND2X1 U1591 ( .A(n1139), .B(n131), .Y(n66) );
  AOI21X1 U1592 ( .A0(n1177), .A1(n133), .B0(n134), .Y(n132) );
  NAND2X1 U1593 ( .A(n522), .B(n534), .Y(n268) );
  NOR2X1 U1594 ( .A(n117), .B(n112), .Y(n110) );
  NAND2X1 U1595 ( .A(n509), .B(n521), .Y(n261) );
  NAND2X1 U1596 ( .A(n535), .B(n545), .Y(n277) );
  CLKINVX1 U1597 ( .A(n346), .Y(n345) );
  CLKINVX1 U1598 ( .A(n328), .Y(n327) );
  CLKINVX1 U1599 ( .A(n326), .Y(n324) );
  CLKINVX1 U1600 ( .A(n344), .Y(n342) );
  OAI21XL U1601 ( .A0(n152), .A1(n144), .B0(n147), .Y(n143) );
  CLKINVX1 U1602 ( .A(n145), .Y(n144) );
  CLKINVX1 U1603 ( .A(n146), .Y(n145) );
  CLKINVX1 U1604 ( .A(n108), .Y(n106) );
  CMPR42X1 U1605 ( .A(n474), .B(n468), .C(n475), .D(n465), .ICI(n471), .S(n462), .ICO(n460), .CO(n461) );
  CMPR42X1 U1606 ( .A(n502), .B(n490), .C(n487), .D(n499), .ICI(n495), .S(n484), .ICO(n482), .CO(n483) );
  NOR2X2 U1607 ( .A(n443), .B(n452), .Y(n213) );
  XNOR2X1 U1608 ( .A(n92), .B(n333), .Y(product[6]) );
  NAND2X1 U1609 ( .A(n1141), .B(n332), .Y(n92) );
  XNOR2X1 U1610 ( .A(n305), .B(n87), .Y(product[11]) );
  NAND2X1 U1611 ( .A(n1142), .B(n350), .Y(n95) );
  CMPR42X1 U1612 ( .A(n547), .B(n541), .C(n548), .D(n538), .ICI(n544), .S(n535), .ICO(n533), .CO(n534) );
  CLKINVX1 U1613 ( .A(n350), .Y(n348) );
  AOI21X1 U1614 ( .A0(n1135), .A1(n302), .B0(n297), .Y(n295) );
  CLKINVX1 U1615 ( .A(n332), .Y(n330) );
  NOR2X2 U1616 ( .A(n592), .B(n597), .Y(n309) );
  NOR2X2 U1617 ( .A(n401), .B(n403), .Y(n139) );
  NAND2X1 U1618 ( .A(n546), .B(n556), .Y(n282) );
  NAND2X1 U1619 ( .A(n435), .B(n442), .Y(n203) );
  XOR2X1 U1620 ( .A(n96), .B(n355), .Y(product[2]) );
  NAND2X1 U1621 ( .A(n1135), .B(n299), .Y(n86) );
  NAND2X1 U1622 ( .A(n336), .B(n339), .Y(n93) );
  NAND2X1 U1623 ( .A(n404), .B(n408), .Y(n147) );
  NAND2X1 U1624 ( .A(n598), .B(n604), .Y(n313) );
  NAND2X1 U1625 ( .A(n803), .B(n787), .Y(n353) );
  NAND2X1 U1626 ( .A(n414), .B(n420), .Y(n165) );
  NAND2X1 U1627 ( .A(n427), .B(n434), .Y(n192) );
  NAND2X1 U1628 ( .A(n413), .B(n409), .Y(n160) );
  NAND2X1 U1629 ( .A(n426), .B(n421), .Y(n179) );
  NAND2X1 U1630 ( .A(n400), .B(n396), .Y(n131) );
  NAND2X1 U1631 ( .A(n401), .B(n403), .Y(n140) );
  NAND2X1 U1632 ( .A(n443), .B(n452), .Y(n214) );
  NAND2X1 U1633 ( .A(n557), .B(n565), .Y(n288) );
  NAND2X1 U1634 ( .A(n621), .B(n785), .Y(n344) );
  CLKINVX1 U1635 ( .A(n338), .Y(n336) );
  CLKINVX1 U1636 ( .A(n431), .Y(n432) );
  CLKINVX1 U1637 ( .A(n469), .Y(n470) );
  NAND2X1 U1638 ( .A(n395), .B(n394), .Y(n122) );
  NAND2X1 U1639 ( .A(n393), .B(n392), .Y(n113) );
  NAND2X1 U1640 ( .A(n391), .B(n634), .Y(n108) );
  CLKINVX1 U1641 ( .A(n391), .Y(n392) );
  CMPR42X1 U1642 ( .A(n661), .B(n705), .C(n481), .D(n491), .ICI(n675), .S(n479), .ICO(n477), .CO(n478) );
  OAI22XL U1643 ( .A0(n851), .A1(n47), .B0(n850), .B1(n46), .Y(n675) );
  OAI22XL U1644 ( .A0(n834), .A1(n52), .B0(n835), .B1(n1013), .Y(n661) );
  OAI22XL U1645 ( .A0(n882), .A1(n34), .B0(n883), .B1(n36), .Y(n705) );
  OR2X1 U1646 ( .A(n771), .B(n678), .Y(n518) );
  AO21X1 U1647 ( .A0(n12), .A1(n9), .B0(n949), .Y(n770) );
  OAI22XL U1648 ( .A0(n866), .A1(n41), .B0(n865), .B1(n40), .Y(n689) );
  OAI22XL U1649 ( .A0(n884), .A1(n34), .B0(n885), .B1(n35), .Y(n707) );
  OAI22XL U1650 ( .A0(n869), .A1(n41), .B0(n868), .B1(n39), .Y(n692) );
  OAI22X1 U1651 ( .A0(n842), .A1(n47), .B0(n841), .B1(n46), .Y(n405) );
  CMPR42X1 U1652 ( .A(n666), .B(n405), .C(n651), .D(n637), .ICI(n402), .S(n401), .ICO(n399), .CO(n400) );
  AO21X1 U1653 ( .A0(n1014), .A1(n46), .B0(n841), .Y(n666) );
  OAI22XL U1654 ( .A0(n808), .A1(n58), .B0(n809), .B1(n60), .Y(n637) );
  OAI22XL U1655 ( .A0(n825), .A1(n54), .B0(n824), .B1(n52), .Y(n651) );
  CMPR42X1 U1656 ( .A(n406), .B(n638), .C(n410), .D(n652), .ICI(n407), .S(n404), .ICO(n402), .CO(n403) );
  OAI22XL U1657 ( .A0(n810), .A1(n60), .B0(n809), .B1(n58), .Y(n638) );
  CLKINVX1 U1658 ( .A(n405), .Y(n406) );
  OAI22XL U1659 ( .A0(n826), .A1(n54), .B0(n825), .B1(n52), .Y(n652) );
  CMPR42X1 U1660 ( .A(n783), .B(n751), .C(n618), .D(n767), .ICI(n799), .S(n615), .ICO(n613), .CO(n614) );
  OAI22XL U1661 ( .A0(n961), .A1(n9), .B0(n962), .B1(n11), .Y(n783) );
  NOR2BX1 U1662 ( .AN(n61), .B(n21), .Y(n751) );
  OAI22XL U1663 ( .A0(n977), .A1(n3), .B0(n978), .B1(n6), .Y(n799) );
  CMPR42X1 U1664 ( .A(n797), .B(n607), .C(n749), .D(n781), .ICI(n608), .S(n605), .ICO(n603), .CO(n604) );
  OAI22XL U1665 ( .A0(n976), .A1(n6), .B0(n975), .B1(n3), .Y(n797) );
  OAI22XL U1666 ( .A0(n928), .A1(n23), .B0(n927), .B1(n21), .Y(n749) );
  OAI22XL U1667 ( .A0(n959), .A1(n9), .B0(n960), .B1(n11), .Y(n781) );
  CMPR42X1 U1668 ( .A(n612), .B(n630), .C(n613), .D(n750), .ICI(n798), .S(n610), .ICO(n608), .CO(n609) );
  OAI22XL U1669 ( .A0(n930), .A1(n22), .B0(n24), .B1(n1038), .Y(n630) );
  OAI22XL U1670 ( .A0(n977), .A1(n1021), .B0(n976), .B1(n3), .Y(n798) );
  OAI22XL U1671 ( .A0(n928), .A1(n21), .B0(n929), .B1(n23), .Y(n750) );
  OAI22XL U1672 ( .A0(n844), .A1(n1014), .B0(n843), .B1(n46), .Y(n668) );
  OAI22XL U1673 ( .A0(n1127), .A1(n60), .B0(n811), .B1(n58), .Y(n640) );
  CMPR42X1 U1674 ( .A(n685), .B(n436), .C(n430), .D(n437), .ICI(n433), .S(n427), .ICO(n425), .CO(n426) );
  CMPR42X1 U1675 ( .A(n702), .B(n454), .C(n455), .D(n446), .ICI(n451), .S(n443), .ICO(n441), .CO(n442) );
  OAI22XL U1676 ( .A0(n880), .A1(n36), .B0(n879), .B1(n34), .Y(n702) );
  OAI22XL U1677 ( .A0(n938), .A1(n18), .B0(n937), .B1(n16), .Y(n759) );
  CMPR42X1 U1678 ( .A(n585), .B(n745), .C(n586), .D(n582), .ICI(n579), .S(n576), .ICO(n574), .CO(n575) );
  OAI22XL U1679 ( .A0(n923), .A1(n21), .B0(n924), .B1(n23), .Y(n745) );
  CMPR42X1 U1680 ( .A(n763), .B(n795), .C(n599), .D(n596), .ICI(n595), .S(n592), .ICO(n590), .CO(n591) );
  OAI22XL U1681 ( .A0(n974), .A1(n6), .B0(n973), .B1(n3), .Y(n795) );
  OAI22XL U1682 ( .A0(n941), .A1(n15), .B0(n942), .B1(n17), .Y(n763) );
  CMPR42X1 U1683 ( .A(n760), .B(n792), .C(n578), .D(n574), .ICI(n569), .S(n566), .ICO(n564), .CO(n565) );
  OAI22XL U1684 ( .A0(n970), .A1(n1031), .B0(n971), .B1(n6), .Y(n792) );
  OAI22XL U1685 ( .A0(n938), .A1(n16), .B0(n939), .B1(n17), .Y(n760) );
  CMPR42X1 U1686 ( .A(n667), .B(n411), .C(n653), .D(n415), .ICI(n412), .S(n409), .ICO(n407), .CO(n408) );
  OAI22XL U1687 ( .A0(n826), .A1(n52), .B0(n827), .B1(n54), .Y(n653) );
  OAI22XL U1688 ( .A0(n843), .A1(n47), .B0(n842), .B1(n46), .Y(n667) );
  OAI22XL U1689 ( .A0(n844), .A1(n46), .B0(n845), .B1(n47), .Y(n669) );
  OAI22XL U1690 ( .A0(n1127), .A1(n58), .B0(n813), .B1(n59), .Y(n641) );
  OAI22XL U1691 ( .A0(n862), .A1(n40), .B0(n863), .B1(n41), .Y(n686) );
  OAI22XL U1692 ( .A0(n815), .A1(n59), .B0(n814), .B1(n57), .Y(n643) );
  NOR2BX1 U1693 ( .AN(n61), .B(n9), .Y(n787) );
  OAI22X1 U1694 ( .A0(n950), .A1(n12), .B0(n949), .B1(n9), .Y(n771) );
  OAI22XL U1695 ( .A0(n820), .A1(n59), .B0(n819), .B1(n57), .Y(n647) );
  OAI22XL U1696 ( .A0(n905), .A1(n30), .B0(n904), .B1(n28), .Y(n726) );
  OAI22XL U1697 ( .A0(n892), .A1(n35), .B0(n891), .B1(n34), .Y(n714) );
  OAI22XL U1698 ( .A0(n958), .A1(n11), .B0(n957), .B1(n9), .Y(n779) );
  CLKINVX1 U1699 ( .A(n397), .Y(n398) );
  OAI22XL U1700 ( .A0(n808), .A1(n60), .B0(n1122), .B1(n58), .Y(n636) );
  OAI22XL U1701 ( .A0(n934), .A1(n16), .B0(n935), .B1(n18), .Y(n756) );
  CMPR42X1 U1702 ( .A(n470), .B(n735), .C(n704), .D(n480), .ICI(n674), .S(n468), .ICO(n466), .CO(n467) );
  OAI22XL U1703 ( .A0(n850), .A1(n47), .B0(n849), .B1(n46), .Y(n674) );
  OAI22XL U1704 ( .A0(n914), .A1(n24), .B0(n913), .B1(n22), .Y(n735) );
  CMPR42X1 U1705 ( .A(n708), .B(n519), .C(n663), .D(n517), .ICI(n526), .S(n515), .ICO(n513), .CO(n514) );
  XNOR2X1 U1706 ( .A(n771), .B(n678), .Y(n519) );
  NAND2X1 U1707 ( .A(n584), .B(n591), .Y(n304) );
  NAND2X1 U1708 ( .A(n576), .B(n583), .Y(n299) );
  OAI22XL U1709 ( .A0(n1130), .A1(n54), .B0(n829), .B1(n52), .Y(n656) );
  CMPR42X1 U1710 ( .A(n469), .B(n734), .C(n645), .D(n688), .ICI(n718), .S(n459), .ICO(n457), .CO(n458) );
  OAI22XL U1711 ( .A0(n864), .A1(n40), .B0(n865), .B1(n41), .Y(n688) );
  CMPR42X1 U1712 ( .A(n697), .B(n727), .C(n570), .D(n791), .ICI(n563), .S(n560), .ICO(n558), .CO(n559) );
  OAI22XL U1713 ( .A0(n970), .A1(n6), .B0(n969), .B1(n1031), .Y(n791) );
  OAI22XL U1714 ( .A0(n874), .A1(n41), .B0(n873), .B1(n39), .Y(n697) );
  CMPR42X1 U1715 ( .A(n747), .B(n716), .C(n601), .D(n779), .ICI(n731), .S(n595), .ICO(n593), .CO(n594) );
  OAI22XL U1716 ( .A0(n910), .A1(n30), .B0(n909), .B1(n28), .Y(n731) );
  OAI22XL U1717 ( .A0(n925), .A1(n21), .B0(n926), .B1(n23), .Y(n747) );
  NOR2BX1 U1718 ( .AN(n61), .B(n34), .Y(n716) );
  CMPR42X1 U1719 ( .A(n736), .B(n690), .C(n720), .D(n488), .ICI(n485), .S(n476), .ICO(n474), .CO(n475) );
  OAI22XL U1720 ( .A0(n894), .A1(n34), .B0(n36), .B1(n1036), .Y(n628) );
  OAI22XL U1721 ( .A0(n1123), .A1(n9), .B0(n957), .B1(n11), .Y(n778) );
  CMPR42X1 U1722 ( .A(n700), .B(n431), .C(n655), .D(n684), .ICI(n428), .S(n424), .ICO(n422), .CO(n423) );
  AO21X1 U1723 ( .A0(n36), .A1(n34), .B0(n877), .Y(n700) );
  OAI22XL U1724 ( .A0(n828), .A1(n52), .B0(n829), .B1(n54), .Y(n655) );
  OAI22XL U1725 ( .A0(n1129), .A1(n24), .B0(n919), .B1(n22), .Y(n741) );
  OAI22XL U1726 ( .A0(n1129), .A1(n22), .B0(n921), .B1(n23), .Y(n742) );
  NAND2X1 U1727 ( .A(n617), .B(n620), .Y(n339) );
  CMPR42X1 U1728 ( .A(n712), .B(n682), .C(n572), .D(n775), .ICI(n743), .S(n563), .ICO(n561), .CO(n562) );
  OAI22XL U1729 ( .A0(n922), .A1(n23), .B0(n921), .B1(n21), .Y(n743) );
  OAI22XL U1730 ( .A0(n889), .A1(n34), .B0(n890), .B1(n35), .Y(n712) );
  OAI22XL U1731 ( .A0(n954), .A1(n12), .B0(n953), .B1(n9), .Y(n775) );
  CLKINVX1 U1732 ( .A(n97), .Y(product[1]) );
  OAI22XL U1733 ( .A0(n1130), .A1(n52), .B0(n831), .B1(n1013), .Y(n657) );
  OAI22XL U1734 ( .A0(n972), .A1(n6), .B0(n971), .B1(n1031), .Y(n793) );
  CMPR42X1 U1735 ( .A(n553), .B(n757), .C(n725), .D(n543), .ICI(n773), .S(n541), .ICO(n539), .CO(n540) );
  OAI22XL U1736 ( .A0(n952), .A1(n12), .B0(n951), .B1(n9), .Y(n773) );
  OAI22XL U1737 ( .A0(n936), .A1(n18), .B0(n935), .B1(n16), .Y(n757) );
  CMPR42X1 U1738 ( .A(n554), .B(n758), .C(n626), .D(n561), .ICI(n774), .S(n552), .ICO(n550), .CO(n551) );
  OAI22XL U1739 ( .A0(n952), .A1(n9), .B0(n953), .B1(n12), .Y(n774) );
  OAI22XL U1740 ( .A0(n870), .A1(n39), .B0(n871), .B1(n41), .Y(n694) );
  ADDFXL U1741 ( .A(n765), .B(n733), .CI(n611), .CO(n606), .S(n607) );
  OAI22XL U1742 ( .A0(n943), .A1(n15), .B0(n944), .B1(n17), .Y(n765) );
  NOR2BX1 U1743 ( .AN(n61), .B(n28), .Y(n733) );
  OAI22XL U1744 ( .A0(n810), .A1(n58), .B0(n811), .B1(n60), .Y(n639) );
  OAI22XL U1745 ( .A0(n871), .A1(n39), .B0(n872), .B1(n41), .Y(n695) );
  ADDFXL U1746 ( .A(n729), .B(n699), .CI(n588), .CO(n580), .S(n581) );
  NOR2BX1 U1747 ( .AN(n61), .B(n39), .Y(n699) );
  ADDFXL U1748 ( .A(n418), .B(n654), .CI(n422), .CO(n415), .S(n416) );
  OAI22XL U1749 ( .A0(n828), .A1(n54), .B0(n827), .B1(n52), .Y(n654) );
  CLKINVX1 U1750 ( .A(n417), .Y(n418) );
  NOR2BX1 U1751 ( .AN(n61), .B(n57), .Y(n649) );
  OR2X1 U1752 ( .A(n788), .B(n679), .Y(n531) );
  NOR2BX1 U1753 ( .AN(n61), .B(n3), .Y(product[0]) );
  OAI22XL U1754 ( .A0(n1122), .A1(n60), .B0(n806), .B1(n58), .Y(n635) );
  XNOR2X1 U1755 ( .A(n990), .B(n25), .Y(n900) );
  XNOR2X1 U1756 ( .A(n995), .B(n43), .Y(n851) );
  XNOR2X1 U1757 ( .A(n995), .B(n37), .Y(n869) );
  XNOR2X1 U1758 ( .A(n995), .B(n31), .Y(n887) );
  XNOR2X1 U1759 ( .A(n996), .B(n43), .Y(n852) );
  XNOR2X1 U1760 ( .A(a[1]), .B(n1), .Y(n982) );
  XNOR2X1 U1761 ( .A(a[1]), .B(n7), .Y(n964) );
  XNOR2X1 U1762 ( .A(a[1]), .B(n13), .Y(n946) );
  XNOR2X1 U1763 ( .A(n990), .B(n37), .Y(n864) );
  XNOR2X1 U1764 ( .A(n990), .B(n31), .Y(n882) );
  XNOR2X1 U1765 ( .A(n990), .B(n19), .Y(n918) );
  XNOR2X1 U1766 ( .A(n990), .B(n13), .Y(n936) );
  XNOR2X1 U1767 ( .A(n988), .B(n7), .Y(n952) );
  XNOR2X1 U1768 ( .A(n990), .B(n7), .Y(n954) );
  XNOR2X1 U1769 ( .A(n995), .B(n25), .Y(n905) );
  XNOR2X1 U1770 ( .A(n988), .B(n1), .Y(n970) );
  XNOR2X1 U1771 ( .A(n995), .B(n19), .Y(n923) );
  XNOR2X1 U1772 ( .A(n990), .B(n1), .Y(n972) );
  XNOR2X1 U1773 ( .A(n995), .B(n13), .Y(n941) );
  XNOR2X1 U1774 ( .A(a[1]), .B(n19), .Y(n928) );
  XNOR2X1 U1775 ( .A(n995), .B(n1), .Y(n977) );
  XNOR2X1 U1776 ( .A(n995), .B(n7), .Y(n959) );
  XNOR2X1 U1777 ( .A(n992), .B(n1), .Y(n974) );
  XNOR2X1 U1778 ( .A(a[1]), .B(n25), .Y(n910) );
  XNOR2X1 U1779 ( .A(a[3]), .B(n55), .Y(n818) );
  XNOR2X1 U1780 ( .A(n986), .B(n31), .Y(n878) );
  XNOR2X1 U1781 ( .A(n997), .B(n55), .Y(n817) );
  XNOR2X1 U1782 ( .A(n997), .B(n43), .Y(n853) );
  XNOR2X1 U1783 ( .A(n996), .B(n55), .Y(n816) );
  XNOR2X1 U1784 ( .A(n996), .B(n49), .Y(n834) );
  XNOR2X1 U1785 ( .A(n986), .B(n43), .Y(n842) );
  XNOR2X1 U1786 ( .A(n997), .B(n37), .Y(n871) );
  XNOR2X1 U1787 ( .A(n997), .B(n25), .Y(n907) );
  XNOR2X1 U1788 ( .A(n996), .B(n37), .Y(n870) );
  XNOR2X1 U1789 ( .A(n987), .B(n7), .Y(n951) );
  XNOR2X1 U1790 ( .A(n997), .B(n31), .Y(n889) );
  XNOR2X1 U1791 ( .A(n996), .B(n19), .Y(n924) );
  XNOR2X1 U1792 ( .A(n996), .B(n13), .Y(n942) );
  XNOR2X1 U1793 ( .A(n997), .B(n13), .Y(n943) );
  XNOR2X1 U1794 ( .A(a[3]), .B(n13), .Y(n944) );
  XNOR2X1 U1795 ( .A(n997), .B(n1), .Y(n979) );
  XNOR2X1 U1796 ( .A(n996), .B(n31), .Y(n888) );
  XNOR2X1 U1797 ( .A(n986), .B(n1), .Y(n968) );
  XNOR2X1 U1798 ( .A(n996), .B(n25), .Y(n906) );
  XNOR2X1 U1799 ( .A(n987), .B(n1), .Y(n969) );
  XNOR2X1 U1800 ( .A(n997), .B(n19), .Y(n925) );
  XNOR2X1 U1801 ( .A(a[3]), .B(n19), .Y(n926) );
  XNOR2X1 U1802 ( .A(n996), .B(n1), .Y(n978) );
  XNOR2X1 U1803 ( .A(n997), .B(n7), .Y(n961) );
  XNOR2X1 U1804 ( .A(n994), .B(n1), .Y(n976) );
  XNOR2X1 U1805 ( .A(n994), .B(n7), .Y(n958) );
  XNOR2X1 U1806 ( .A(a[2]), .B(n1), .Y(n981) );
  XNOR2X1 U1807 ( .A(n989), .B(n19), .Y(n917) );
  XNOR2X1 U1808 ( .A(a[2]), .B(n31), .Y(n891) );
  XNOR2X1 U1809 ( .A(a[2]), .B(n49), .Y(n837) );
  XNOR2X1 U1810 ( .A(n993), .B(n13), .Y(n939) );
  XNOR2X1 U1811 ( .A(n991), .B(n7), .Y(n955) );
  XNOR2X1 U1812 ( .A(a[2]), .B(n7), .Y(n963) );
  XNOR2X1 U1813 ( .A(n989), .B(n13), .Y(n935) );
  XNOR2X1 U1814 ( .A(a[2]), .B(n43), .Y(n855) );
  XNOR2X1 U1815 ( .A(n991), .B(n19), .Y(n919) );
  XNOR2X1 U1816 ( .A(a[2]), .B(n37), .Y(n873) );
  XNOR2X1 U1817 ( .A(a[2]), .B(n25), .Y(n909) );
  XNOR2X1 U1818 ( .A(n993), .B(n7), .Y(n957) );
  XNOR2X1 U1819 ( .A(a[2]), .B(n19), .Y(n927) );
  XNOR2X1 U1820 ( .A(n993), .B(n1), .Y(n975) );
  XNOR2X1 U1821 ( .A(n985), .B(n25), .Y(n895) );
  XNOR2X1 U1822 ( .A(n985), .B(n31), .Y(n877) );
  XNOR2X1 U1823 ( .A(n985), .B(n1), .Y(n967) );
  CLKINVX1 U1824 ( .A(n13), .Y(n1039) );
  CMPR42X1 U1825 ( .A(n580), .B(n698), .C(n744), .D(n571), .ICI(n577), .S(n569), .ICO(n567), .CO(n568) );
  OAI22XL U1826 ( .A0(n874), .A1(n39), .B0(n875), .B1(n41), .Y(n698) );
  OAI22XL U1827 ( .A0(n923), .A1(n23), .B0(n922), .B1(n21), .Y(n744) );
  XNOR2X1 U1828 ( .A(n61), .B(n37), .Y(n875) );
  CMPR42X1 U1829 ( .A(n715), .B(n762), .C(n594), .D(n590), .ICI(n587), .S(n584), .ICO(n582), .CO(n583) );
  OAI22XL U1830 ( .A0(n892), .A1(n1026), .B0(n893), .B1(n35), .Y(n715) );
  OAI22XL U1831 ( .A0(n941), .A1(n17), .B0(n940), .B1(n15), .Y(n762) );
  XNOR2X1 U1832 ( .A(n61), .B(n31), .Y(n893) );
  CLKBUFX3 U1833 ( .A(n1020), .Y(n12) );
  CLKINVX1 U1834 ( .A(n7), .Y(n1040) );
  OAI22XL U1835 ( .A0(n876), .A1(n40), .B0(n41), .B1(n1035), .Y(n627) );
  CLKINVX1 U1836 ( .A(n37), .Y(n1035) );
  OAI22XL U1837 ( .A0(n912), .A1(n28), .B0(n30), .B1(n1037), .Y(n629) );
  CLKINVX1 U1838 ( .A(n25), .Y(n1037) );
  XNOR2X1 U1839 ( .A(n986), .B(n55), .Y(n806) );
  CLKBUFX3 U1840 ( .A(n1023), .Y(n52) );
  CLKBUFX3 U1841 ( .A(n1022), .Y(n58) );
  CLKBUFX3 U1842 ( .A(n1024), .Y(n46) );
  CLKBUFX3 U1843 ( .A(n1025), .Y(n40) );
  CLKBUFX3 U1844 ( .A(n1022), .Y(n57) );
  CLKBUFX3 U1845 ( .A(n1025), .Y(n39) );
  CLKBUFX3 U1846 ( .A(n1029), .Y(n15) );
  CLKBUFX3 U1847 ( .A(n1028), .Y(n21) );
  CLKBUFX3 U1848 ( .A(n1012), .Y(n59) );
  CLKBUFX3 U1849 ( .A(n1016), .Y(n35) );
  CLKBUFX3 U1850 ( .A(n1018), .Y(n23) );
  CLKBUFX3 U1851 ( .A(n1013), .Y(n54) );
  CLKBUFX3 U1852 ( .A(n1012), .Y(n60) );
  CLKBUFX3 U1853 ( .A(n1016), .Y(n36) );
  CLKINVX1 U1854 ( .A(n31), .Y(n1036) );
  CLKINVX1 U1855 ( .A(n19), .Y(n1038) );
  CLKINVX1 U1856 ( .A(n55), .Y(n1032) );
  XNOR2X1 U1857 ( .A(n985), .B(n55), .Y(n805) );
  XOR2X1 U1858 ( .A(n1133), .B(b[19]), .Y(n1002) );
  NAND2X1 U1859 ( .A(n1007), .B(n1027), .Y(n1017) );
  XOR2X1 U1860 ( .A(b[8]), .B(b[9]), .Y(n1007) );
  XOR2X1 U1861 ( .A(b[14]), .B(b[15]), .Y(n1004) );
  NAND2X1 U1862 ( .A(n1005), .B(n1025), .Y(n1015) );
  XOR2X1 U1863 ( .A(b[12]), .B(b[13]), .Y(n1005) );
  XOR2X1 U1864 ( .A(b[4]), .B(b[5]), .Y(n1009) );
endmodule


module CONV_DW01_add_5 ( A, B, CI, SUM, CO );
  input [43:0] A;
  input [43:0] B;
  output [43:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n47, n48, n53, n54, n55, n56, n57, n59, n61, n62, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n124, n125, n127, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n149, n150, n151, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n166, n168, n171, n173, n174, n175, n176,
         n177, n178, n179, n181, n183, n184, n185, n186, n187, n188, n190,
         n192, n193, n194, n195, n196, n197, n198, n199, n201, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n249, n251,
         n254, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n271, n273, n276, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n306, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n321, n324, n325, n326, n328, n330, n332, n333,
         n334, n340, n341, n342, n343, n344, n345, n346, n347, n350, n351,
         n354, n355, n356, n357, n358, n359, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517;

  INVX1 U411 ( .A(n93), .Y(n91) );
  NOR2X2 U412 ( .A(B[6]), .B(A[6]), .Y(n295) );
  NAND2XL U413 ( .A(n65), .B(n68), .Y(n5) );
  INVX1 U414 ( .A(n68), .Y(n66) );
  OAI21X4 U415 ( .A0(n312), .A1(n310), .B0(n311), .Y(n309) );
  AOI21X4 U416 ( .A0(n313), .A1(n317), .B0(n314), .Y(n312) );
  OAI21X2 U417 ( .A0(n228), .A1(n234), .B0(n229), .Y(n227) );
  AOI21X1 U418 ( .A0(n227), .A1(n218), .B0(n219), .Y(n217) );
  NAND2X2 U419 ( .A(B[10]), .B(A[10]), .Y(n278) );
  NAND2X2 U420 ( .A(B[21]), .B(A[21]), .Y(n221) );
  CLKINVX1 U421 ( .A(n198), .Y(n196) );
  NAND2X1 U422 ( .A(B[0]), .B(A[0]), .Y(n319) );
  NOR2X1 U423 ( .A(n223), .B(n220), .Y(n218) );
  NOR2X1 U424 ( .A(n102), .B(n95), .Y(n93) );
  NOR2X1 U425 ( .A(n228), .B(n233), .Y(n226) );
  CLKINVX1 U426 ( .A(n168), .Y(n166) );
  OAI21X1 U427 ( .A0(n239), .A1(n243), .B0(n240), .Y(n238) );
  NOR2X1 U428 ( .A(n242), .B(n239), .Y(n237) );
  OA21XL U429 ( .A0(n95), .A1(n103), .B0(n96), .Y(n510) );
  AOI21X1 U430 ( .A0(n281), .A1(n289), .B0(n282), .Y(n280) );
  OAI21X1 U431 ( .A0(n292), .A1(n290), .B0(n291), .Y(n289) );
  OAI21XL U432 ( .A0(n75), .A1(n85), .B0(n76), .Y(n74) );
  NOR2X1 U433 ( .A(n71), .B(n109), .Y(n69) );
  NAND2X1 U434 ( .A(B[14]), .B(A[14]), .Y(n256) );
  OR2X1 U435 ( .A(B[24]), .B(A[24]), .Y(n502) );
  OAI21X2 U436 ( .A0(n209), .A1(n213), .B0(n210), .Y(n208) );
  NAND2X1 U437 ( .A(B[28]), .B(A[28]), .Y(n168) );
  OAI21XL U438 ( .A0(n155), .A1(n147), .B0(n150), .Y(n146) );
  INVX3 U439 ( .A(n175), .Y(n174) );
  NOR2X1 U440 ( .A(B[19]), .B(A[19]), .Y(n228) );
  NAND2X1 U441 ( .A(B[5]), .B(A[5]), .Y(n299) );
  XNOR2X1 U442 ( .A(n55), .B(n3), .Y(SUM[42]) );
  OAI21X1 U443 ( .A0(n136), .A1(n127), .B0(n124), .Y(n122) );
  XOR2X1 U444 ( .A(n225), .B(n25), .Y(SUM[20]) );
  OAI21XL U445 ( .A0(n214), .A1(n506), .B0(n213), .Y(n211) );
  OAI21XL U446 ( .A0(n214), .A1(n194), .B0(n195), .Y(n193) );
  XNOR2X1 U447 ( .A(n133), .B(n12), .Y(SUM[33]) );
  OAI21X1 U448 ( .A0(n136), .A1(n116), .B0(n117), .Y(n115) );
  XNOR2X1 U449 ( .A(n86), .B(n7), .Y(SUM[38]) );
  XNOR2X1 U450 ( .A(n97), .B(n8), .Y(SUM[37]) );
  XNOR2X1 U451 ( .A(n104), .B(n9), .Y(SUM[36]) );
  CLKINVX1 U452 ( .A(n315), .Y(n313) );
  XNOR2X1 U453 ( .A(n48), .B(n2), .Y(SUM[43]) );
  NAND2X1 U454 ( .A(B[11]), .B(A[11]), .Y(n273) );
  OR2X2 U455 ( .A(B[28]), .B(A[28]), .Y(n495) );
  OR2XL U456 ( .A(B[36]), .B(A[41]), .Y(n496) );
  OR2X1 U457 ( .A(B[11]), .B(A[11]), .Y(n497) );
  OR2X1 U458 ( .A(B[14]), .B(A[14]), .Y(n498) );
  OR2X1 U459 ( .A(B[26]), .B(A[26]), .Y(n499) );
  OR2X1 U460 ( .A(B[27]), .B(A[27]), .Y(n500) );
  OR2X1 U461 ( .A(B[10]), .B(A[10]), .Y(n501) );
  INVX1 U462 ( .A(n67), .Y(n65) );
  OR2X1 U463 ( .A(B[3]), .B(A[3]), .Y(n503) );
  OR2X8 U464 ( .A(B[15]), .B(A[15]), .Y(n504) );
  OR2X1 U465 ( .A(B[25]), .B(A[25]), .Y(n505) );
  NAND2X1 U466 ( .A(B[34]), .B(A[34]), .Y(n121) );
  CLKINVX1 U467 ( .A(n110), .Y(n108) );
  CLKBUFX3 U468 ( .A(n120), .Y(n507) );
  CLKINVX1 U469 ( .A(n507), .Y(n118) );
  NOR2X1 U470 ( .A(B[36]), .B(A[36]), .Y(n102) );
  OAI21X1 U471 ( .A0(n220), .A1(n224), .B0(n221), .Y(n219) );
  NOR2X6 U472 ( .A(n514), .B(n70), .Y(n1) );
  NOR2X1 U473 ( .A(B[34]), .B(A[34]), .Y(n120) );
  INVX1 U474 ( .A(n215), .Y(n214) );
  AO21XL U475 ( .A0(n174), .A1(n500), .B0(n171), .Y(n511) );
  XNOR2XL U476 ( .A(n174), .B(n18), .Y(SUM[27]) );
  OAI21X1 U477 ( .A0(n136), .A1(n134), .B0(n135), .Y(n133) );
  INVX3 U478 ( .A(n137), .Y(n136) );
  NAND2XL U479 ( .A(n346), .B(n240), .Y(n28) );
  NAND2X1 U480 ( .A(B[17]), .B(A[17]), .Y(n240) );
  AOI21X4 U481 ( .A0(n267), .A1(n259), .B0(n260), .Y(n258) );
  OAI21X1 U482 ( .A0(n261), .A1(n265), .B0(n262), .Y(n260) );
  OAI21X1 U483 ( .A0(n136), .A1(n109), .B0(n106), .Y(n104) );
  NAND2X2 U484 ( .A(B[22]), .B(A[22]), .Y(n213) );
  OAI21X1 U485 ( .A0(n136), .A1(n87), .B0(n88), .Y(n86) );
  XOR2X1 U486 ( .A(n1), .B(n5), .Y(SUM[40]) );
  NOR2X4 U487 ( .A(B[9]), .B(A[9]), .Y(n283) );
  NAND2X2 U488 ( .A(B[9]), .B(A[9]), .Y(n284) );
  OAI21X1 U489 ( .A0(n136), .A1(n98), .B0(n99), .Y(n97) );
  INVXL U490 ( .A(n242), .Y(n347) );
  NOR2X4 U491 ( .A(B[16]), .B(A[16]), .Y(n242) );
  BUFX8 U492 ( .A(n212), .Y(n506) );
  NAND2X4 U493 ( .A(B[15]), .B(A[15]), .Y(n251) );
  OAI21X1 U494 ( .A0(n1), .A1(n516), .B0(n515), .Y(n48) );
  OAI21X1 U495 ( .A0(n1), .A1(n56), .B0(n57), .Y(n55) );
  XNOR2X4 U496 ( .A(n62), .B(n4), .Y(SUM[41]) );
  OAI21X1 U497 ( .A0(n1), .A1(n67), .B0(n68), .Y(n62) );
  INVXL U498 ( .A(n149), .Y(n333) );
  NOR2X2 U499 ( .A(n149), .B(n142), .Y(n140) );
  NOR2X2 U500 ( .A(n113), .B(n507), .Y(n111) );
  INVXL U501 ( .A(n223), .Y(n343) );
  OAI21X2 U502 ( .A0(n225), .A1(n223), .B0(n224), .Y(n222) );
  NOR2X2 U503 ( .A(B[20]), .B(A[20]), .Y(n223) );
  AND2X4 U504 ( .A(n235), .B(n226), .Y(n508) );
  NOR2X6 U505 ( .A(n508), .B(n227), .Y(n225) );
  INVXL U506 ( .A(n236), .Y(n235) );
  NAND2X2 U507 ( .A(B[31]), .B(A[31]), .Y(n143) );
  NOR2X6 U508 ( .A(B[31]), .B(A[31]), .Y(n142) );
  AOI21X2 U509 ( .A0(n130), .A1(n111), .B0(n112), .Y(n110) );
  OAI21X1 U510 ( .A0(n304), .A1(n302), .B0(n303), .Y(n301) );
  OR2XL U511 ( .A(B[32]), .B(A[32]), .Y(n509) );
  NAND2X2 U512 ( .A(B[25]), .B(A[25]), .Y(n192) );
  NOR2X6 U513 ( .A(B[12]), .B(A[12]), .Y(n264) );
  NAND2X6 U514 ( .A(B[12]), .B(A[12]), .Y(n265) );
  NAND2X2 U515 ( .A(B[36]), .B(A[36]), .Y(n103) );
  NOR2X6 U516 ( .A(B[21]), .B(A[21]), .Y(n220) );
  INVX1 U517 ( .A(n155), .Y(n153) );
  INVXL U518 ( .A(n207), .Y(n205) );
  NAND2X1 U519 ( .A(n328), .B(n114), .Y(n10) );
  NAND2X1 U520 ( .A(B[35]), .B(A[35]), .Y(n114) );
  NAND2X4 U521 ( .A(B[32]), .B(A[32]), .Y(n135) );
  NAND2X4 U522 ( .A(B[16]), .B(A[16]), .Y(n243) );
  NAND2X4 U523 ( .A(B[30]), .B(A[30]), .Y(n150) );
  NAND2X4 U524 ( .A(B[20]), .B(A[20]), .Y(n224) );
  NOR2X1 U525 ( .A(B[30]), .B(A[30]), .Y(n149) );
  NOR2X1 U526 ( .A(B[32]), .B(A[32]), .Y(n134) );
  NAND2X1 U527 ( .A(B[2]), .B(A[2]), .Y(n311) );
  NAND2X1 U528 ( .A(n207), .B(n502), .Y(n198) );
  INVXL U529 ( .A(n113), .Y(n328) );
  OAI21X1 U530 ( .A0(n113), .A1(n121), .B0(n114), .Y(n112) );
  NOR2X2 U531 ( .A(n506), .B(n209), .Y(n207) );
  NOR2X2 U532 ( .A(B[8]), .B(A[8]), .Y(n286) );
  NOR2X2 U533 ( .A(n198), .B(n178), .Y(n176) );
  NOR2X1 U534 ( .A(B[22]), .B(A[22]), .Y(n212) );
  NAND2X2 U535 ( .A(B[8]), .B(A[8]), .Y(n287) );
  NAND2X1 U536 ( .A(n65), .B(n496), .Y(n56) );
  AOI21X1 U537 ( .A0(n94), .A1(n73), .B0(n74), .Y(n72) );
  AOI21X2 U538 ( .A0(n237), .A1(n245), .B0(n238), .Y(n236) );
  NOR2X2 U539 ( .A(B[2]), .B(A[2]), .Y(n310) );
  NOR2X1 U540 ( .A(B[5]), .B(A[5]), .Y(n298) );
  NAND2X1 U541 ( .A(B[3]), .B(A[3]), .Y(n308) );
  NAND2XL U542 ( .A(B[4]), .B(A[4]), .Y(n303) );
  NAND2X1 U543 ( .A(B[1]), .B(A[1]), .Y(n316) );
  NAND2X1 U544 ( .A(B[7]), .B(A[7]), .Y(n291) );
  AND2X2 U545 ( .A(n137), .B(n69), .Y(n514) );
  OAI21X1 U546 ( .A0(n110), .A1(n71), .B0(n72), .Y(n70) );
  NOR2X1 U547 ( .A(n131), .B(n134), .Y(n129) );
  AOI21X2 U548 ( .A0(n495), .A1(n171), .B0(n166), .Y(n164) );
  NOR2X1 U549 ( .A(n283), .B(n286), .Y(n281) );
  OAI21X2 U550 ( .A0(n258), .A1(n246), .B0(n247), .Y(n245) );
  NOR2X1 U551 ( .A(B[18]), .B(A[18]), .Y(n233) );
  NOR2X1 U552 ( .A(B[1]), .B(A[1]), .Y(n315) );
  NOR2X1 U553 ( .A(B[7]), .B(A[7]), .Y(n290) );
  NOR2X1 U554 ( .A(B[4]), .B(A[4]), .Y(n302) );
  CLKINVX1 U555 ( .A(n129), .Y(n127) );
  INVXL U556 ( .A(n53), .Y(n321) );
  AOI21X1 U557 ( .A0(n108), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U558 ( .A0(n309), .A1(n503), .B0(n306), .Y(n304) );
  NAND2X1 U559 ( .A(B[26]), .B(A[26]), .Y(n183) );
  NAND2X1 U560 ( .A(B[13]), .B(A[13]), .Y(n262) );
  NOR2X2 U561 ( .A(B[29]), .B(A[29]), .Y(n158) );
  NAND2X2 U562 ( .A(B[18]), .B(A[18]), .Y(n234) );
  NAND2X1 U563 ( .A(B[6]), .B(A[6]), .Y(n296) );
  NAND2X2 U564 ( .A(n129), .B(n111), .Y(n109) );
  INVXL U565 ( .A(n510), .Y(n90) );
  NAND2XL U566 ( .A(n80), .B(n107), .Y(n78) );
  INVXL U567 ( .A(n130), .Y(n124) );
  AOI21X2 U568 ( .A0(n215), .A1(n176), .B0(n177), .Y(n175) );
  OAI21X2 U569 ( .A0(n199), .A1(n178), .B0(n179), .Y(n177) );
  NAND2X2 U570 ( .A(n495), .B(n500), .Y(n163) );
  INVXL U571 ( .A(n199), .Y(n197) );
  AOI21XL U572 ( .A0(n197), .A1(n187), .B0(n190), .Y(n186) );
  OAI21X4 U573 ( .A0(n216), .A1(n236), .B0(n217), .Y(n215) );
  NAND2X2 U574 ( .A(n218), .B(n226), .Y(n216) );
  OAI21X2 U575 ( .A0(n164), .A1(n158), .B0(n159), .Y(n157) );
  NAND2XL U576 ( .A(n324), .B(n76), .Y(n6) );
  OAI21X1 U577 ( .A0(n136), .A1(n78), .B0(n79), .Y(n77) );
  INVXL U578 ( .A(n75), .Y(n324) );
  NAND2XL U579 ( .A(n325), .B(n85), .Y(n7) );
  INVXL U580 ( .A(n84), .Y(n325) );
  OAI21X1 U581 ( .A0(n283), .A1(n287), .B0(n284), .Y(n282) );
  OAI21XL U582 ( .A0(n95), .A1(n103), .B0(n96), .Y(n94) );
  OAI21X2 U583 ( .A0(n131), .A1(n135), .B0(n132), .Y(n130) );
  OAI21X2 U584 ( .A0(n280), .A1(n268), .B0(n269), .Y(n267) );
  NAND2X2 U585 ( .A(n497), .B(n501), .Y(n268) );
  NAND2X2 U586 ( .A(n504), .B(n498), .Y(n246) );
  NOR2X4 U587 ( .A(n158), .B(n163), .Y(n156) );
  AOI21X2 U588 ( .A0(n496), .A1(n66), .B0(n59), .Y(n57) );
  XOR2XL U589 ( .A(n136), .B(n13), .Y(SUM[32]) );
  NAND2XL U590 ( .A(n334), .B(n159), .Y(n16) );
  XNOR2X1 U591 ( .A(n511), .B(n17), .Y(SUM[28]) );
  NAND2XL U592 ( .A(n502), .B(n203), .Y(n21) );
  NAND2XL U593 ( .A(n340), .B(n210), .Y(n22) );
  INVXL U594 ( .A(n209), .Y(n340) );
  XOR2XL U595 ( .A(n214), .B(n23), .Y(SUM[22]) );
  NAND2XL U596 ( .A(n341), .B(n213), .Y(n23) );
  NAND2XL U597 ( .A(n344), .B(n229), .Y(n26) );
  AOI21XL U598 ( .A0(n235), .A1(n345), .B0(n232), .Y(n230) );
  INVXL U599 ( .A(n228), .Y(n344) );
  INVXL U600 ( .A(n102), .Y(n100) );
  XOR2XL U601 ( .A(n244), .B(n29), .Y(SUM[16]) );
  XNOR2X1 U602 ( .A(n512), .B(n30), .Y(SUM[15]) );
  AO21XL U603 ( .A0(n257), .A1(n498), .B0(n254), .Y(n512) );
  XNOR2XL U604 ( .A(n235), .B(n27), .Y(SUM[18]) );
  XOR2XL U605 ( .A(n266), .B(n33), .Y(SUM[12]) );
  XNOR2X1 U606 ( .A(n513), .B(n34), .Y(SUM[11]) );
  AO21XL U607 ( .A0(n279), .A1(n501), .B0(n276), .Y(n513) );
  XNOR2XL U608 ( .A(n257), .B(n31), .Y(SUM[14]) );
  XOR2XL U609 ( .A(n288), .B(n37), .Y(SUM[8]) );
  XOR2XL U610 ( .A(n292), .B(n38), .Y(SUM[7]) );
  INVXL U611 ( .A(n295), .Y(n357) );
  XNOR2XL U612 ( .A(n279), .B(n35), .Y(SUM[10]) );
  XOR2XL U613 ( .A(n304), .B(n41), .Y(SUM[4]) );
  XNOR2XL U614 ( .A(n309), .B(n42), .Y(SUM[3]) );
  NAND2X2 U615 ( .A(B[27]), .B(A[27]), .Y(n173) );
  NAND2XL U616 ( .A(B[36]), .B(A[43]), .Y(n47) );
  NAND2XL U617 ( .A(B[36]), .B(A[40]), .Y(n68) );
  NOR2X4 U618 ( .A(B[35]), .B(A[35]), .Y(n113) );
  NOR2X1 U619 ( .A(B[36]), .B(A[42]), .Y(n53) );
  NAND2XL U620 ( .A(B[36]), .B(A[41]), .Y(n61) );
  NAND2XL U621 ( .A(B[36]), .B(A[42]), .Y(n54) );
  NOR2XL U622 ( .A(B[36]), .B(A[40]), .Y(n67) );
  OR2XL U623 ( .A(B[36]), .B(A[43]), .Y(n517) );
  XOR2XL U624 ( .A(n43), .B(n312), .Y(SUM[2]) );
  XNOR2XL U625 ( .A(n44), .B(n317), .Y(SUM[1]) );
  NOR2XL U626 ( .A(B[0]), .B(A[0]), .Y(n318) );
  NAND2BXL U627 ( .AN(n318), .B(n319), .Y(n45) );
  OAI21X4 U628 ( .A0(n175), .A1(n138), .B0(n139), .Y(n137) );
  NAND2X1 U629 ( .A(n107), .B(n89), .Y(n87) );
  CLKINVX1 U630 ( .A(n196), .Y(n194) );
  CLKINVX1 U631 ( .A(n109), .Y(n107) );
  AOI21X1 U632 ( .A0(n108), .A1(n89), .B0(n90), .Y(n88) );
  CLKINVX1 U633 ( .A(n91), .Y(n89) );
  CLKINVX1 U634 ( .A(n108), .Y(n106) );
  NAND2X1 U635 ( .A(n196), .B(n187), .Y(n185) );
  CLKINVX1 U636 ( .A(n163), .Y(n161) );
  CLKINVX1 U637 ( .A(n197), .Y(n195) );
  NAND2X1 U638 ( .A(n93), .B(n73), .Y(n71) );
  NAND2X1 U639 ( .A(n499), .B(n505), .Y(n178) );
  NOR2X1 U640 ( .A(n91), .B(n84), .Y(n80) );
  CLKINVX1 U641 ( .A(n156), .Y(n154) );
  CLKINVX1 U642 ( .A(n157), .Y(n155) );
  CLKINVX1 U643 ( .A(n127), .Y(n125) );
  NOR2X1 U644 ( .A(n154), .B(n147), .Y(n145) );
  CLKINVX1 U645 ( .A(n164), .Y(n162) );
  NAND2X1 U646 ( .A(n107), .B(n100), .Y(n98) );
  NAND2X1 U647 ( .A(n125), .B(n118), .Y(n116) );
  CLKINVX1 U648 ( .A(n267), .Y(n266) );
  CLKINVX1 U649 ( .A(n245), .Y(n244) );
  CLKINVX1 U650 ( .A(n258), .Y(n257) );
  CLKINVX1 U651 ( .A(n208), .Y(n206) );
  CLKINVX1 U652 ( .A(n188), .Y(n187) );
  CLKINVX1 U653 ( .A(n505), .Y(n188) );
  CLKINVX1 U654 ( .A(n289), .Y(n288) );
  CLKINVX1 U655 ( .A(n280), .Y(n279) );
  CLKINVX1 U656 ( .A(n301), .Y(n300) );
  NAND2X1 U657 ( .A(n496), .B(n61), .Y(n4) );
  NAND2X1 U658 ( .A(n321), .B(n54), .Y(n3) );
  NOR2X1 U659 ( .A(n84), .B(n75), .Y(n73) );
  NOR2X1 U660 ( .A(n264), .B(n261), .Y(n259) );
  AOI21X1 U661 ( .A0(n208), .A1(n502), .B0(n201), .Y(n199) );
  CLKINVX1 U662 ( .A(n203), .Y(n201) );
  AOI21X1 U663 ( .A0(n497), .A1(n276), .B0(n271), .Y(n269) );
  CLKINVX1 U664 ( .A(n273), .Y(n271) );
  NAND2X1 U665 ( .A(n140), .B(n156), .Y(n138) );
  AOI21X1 U666 ( .A0(n157), .A1(n140), .B0(n141), .Y(n139) );
  AOI21X1 U667 ( .A0(n504), .A1(n254), .B0(n249), .Y(n247) );
  CLKINVX1 U668 ( .A(n308), .Y(n306) );
  AOI21X1 U669 ( .A0(n293), .A1(n301), .B0(n294), .Y(n292) );
  NOR2X1 U670 ( .A(n295), .B(n298), .Y(n293) );
  OAI21XL U671 ( .A0(n295), .A1(n299), .B0(n296), .Y(n294) );
  CLKINVX1 U672 ( .A(n316), .Y(n314) );
  CLKINVX1 U673 ( .A(n61), .Y(n59) );
  NAND2X1 U674 ( .A(n100), .B(n103), .Y(n9) );
  XNOR2X1 U675 ( .A(n77), .B(n6), .Y(SUM[39]) );
  NAND2X1 U676 ( .A(n326), .B(n96), .Y(n8) );
  CLKINVX1 U677 ( .A(n95), .Y(n326) );
  XNOR2X1 U678 ( .A(n122), .B(n11), .Y(SUM[34]) );
  NAND2X1 U679 ( .A(n118), .B(n121), .Y(n11) );
  NAND2X1 U680 ( .A(n500), .B(n173), .Y(n18) );
  XNOR2X1 U681 ( .A(n211), .B(n22), .Y(SUM[23]) );
  NAND2X1 U682 ( .A(n330), .B(n132), .Y(n12) );
  CLKINVX1 U683 ( .A(n131), .Y(n330) );
  XNOR2X1 U684 ( .A(n115), .B(n10), .Y(SUM[35]) );
  OAI21XL U685 ( .A0(n142), .A1(n150), .B0(n143), .Y(n141) );
  AOI21X1 U686 ( .A0(n80), .A1(n108), .B0(n81), .Y(n79) );
  OAI21XL U687 ( .A0(n510), .A1(n84), .B0(n85), .Y(n81) );
  CLKINVX1 U688 ( .A(n103), .Y(n101) );
  AOI21X1 U689 ( .A0(n130), .A1(n118), .B0(n119), .Y(n117) );
  CLKINVX1 U690 ( .A(n121), .Y(n119) );
  AOI21X1 U691 ( .A0(n499), .A1(n190), .B0(n181), .Y(n179) );
  CLKINVX1 U692 ( .A(n183), .Y(n181) );
  XNOR2X1 U693 ( .A(n184), .B(n19), .Y(SUM[26]) );
  NAND2X1 U694 ( .A(n499), .B(n183), .Y(n19) );
  OAI21XL U695 ( .A0(n214), .A1(n185), .B0(n186), .Y(n184) );
  XNOR2X1 U696 ( .A(n193), .B(n20), .Y(SUM[25]) );
  NAND2X1 U697 ( .A(n187), .B(n192), .Y(n20) );
  XNOR2X1 U698 ( .A(n204), .B(n21), .Y(SUM[24]) );
  OAI21XL U699 ( .A0(n214), .A1(n205), .B0(n206), .Y(n204) );
  CLKINVX1 U700 ( .A(n333), .Y(n147) );
  CLKINVX1 U701 ( .A(n192), .Y(n190) );
  CLKINVX1 U702 ( .A(n173), .Y(n171) );
  CLKINVX1 U703 ( .A(n256), .Y(n254) );
  CLKINVX1 U704 ( .A(n278), .Y(n276) );
  XOR2X1 U705 ( .A(n144), .B(n14), .Y(SUM[31]) );
  NAND2X1 U706 ( .A(n332), .B(n143), .Y(n14) );
  AOI21X1 U707 ( .A0(n174), .A1(n145), .B0(n146), .Y(n144) );
  CLKINVX1 U708 ( .A(n142), .Y(n332) );
  XOR2X1 U709 ( .A(n151), .B(n15), .Y(SUM[30]) );
  NAND2X1 U710 ( .A(n333), .B(n150), .Y(n15) );
  AOI21X1 U711 ( .A0(n174), .A1(n156), .B0(n153), .Y(n151) );
  XOR2X1 U712 ( .A(n160), .B(n16), .Y(SUM[29]) );
  AOI21X1 U713 ( .A0(n174), .A1(n161), .B0(n162), .Y(n160) );
  CLKINVX1 U714 ( .A(n158), .Y(n334) );
  NAND2X1 U715 ( .A(n495), .B(n168), .Y(n17) );
  NAND2X1 U716 ( .A(n509), .B(n135), .Y(n13) );
  CLKINVX1 U717 ( .A(n251), .Y(n249) );
  OA21XL U718 ( .A0(n57), .A1(n53), .B0(n54), .Y(n515) );
  OR2X1 U719 ( .A(n56), .B(n53), .Y(n516) );
  XNOR2X1 U720 ( .A(n222), .B(n24), .Y(SUM[21]) );
  NAND2X1 U721 ( .A(n342), .B(n221), .Y(n24) );
  CLKINVX1 U722 ( .A(n220), .Y(n342) );
  NAND2X1 U723 ( .A(n498), .B(n256), .Y(n31) );
  NAND2X1 U724 ( .A(n345), .B(n234), .Y(n27) );
  CLKINVX1 U725 ( .A(n233), .Y(n345) );
  XNOR2X1 U726 ( .A(n241), .B(n28), .Y(SUM[17]) );
  OAI21XL U727 ( .A0(n244), .A1(n242), .B0(n243), .Y(n241) );
  CLKINVX1 U728 ( .A(n239), .Y(n346) );
  XNOR2X1 U729 ( .A(n263), .B(n32), .Y(SUM[13]) );
  NAND2X1 U730 ( .A(n350), .B(n262), .Y(n32) );
  OAI21XL U731 ( .A0(n266), .A1(n264), .B0(n265), .Y(n263) );
  CLKINVX1 U732 ( .A(n261), .Y(n350) );
  CLKINVX1 U733 ( .A(n319), .Y(n317) );
  NAND2X1 U734 ( .A(n347), .B(n243), .Y(n29) );
  XOR2X1 U735 ( .A(n230), .B(n26), .Y(SUM[19]) );
  NAND2X1 U736 ( .A(n504), .B(n251), .Y(n30) );
  CLKINVX1 U737 ( .A(n506), .Y(n341) );
  NAND2X1 U738 ( .A(n343), .B(n224), .Y(n25) );
  CLKINVX1 U739 ( .A(n234), .Y(n232) );
  NAND2X1 U740 ( .A(n501), .B(n278), .Y(n35) );
  XNOR2X1 U741 ( .A(n285), .B(n36), .Y(SUM[9]) );
  NAND2X1 U742 ( .A(n354), .B(n284), .Y(n36) );
  OAI21XL U743 ( .A0(n288), .A1(n286), .B0(n287), .Y(n285) );
  CLKINVX1 U744 ( .A(n283), .Y(n354) );
  NAND2X1 U745 ( .A(n351), .B(n265), .Y(n33) );
  CLKINVX1 U746 ( .A(n264), .Y(n351) );
  NAND2X1 U747 ( .A(n355), .B(n287), .Y(n37) );
  CLKINVX1 U748 ( .A(n286), .Y(n355) );
  NAND2X1 U749 ( .A(n497), .B(n273), .Y(n34) );
  NAND2X1 U750 ( .A(n356), .B(n291), .Y(n38) );
  CLKINVX1 U751 ( .A(n290), .Y(n356) );
  XNOR2X1 U752 ( .A(n297), .B(n39), .Y(SUM[6]) );
  NAND2X1 U753 ( .A(n357), .B(n296), .Y(n39) );
  OAI21XL U754 ( .A0(n300), .A1(n298), .B0(n299), .Y(n297) );
  NAND2X1 U755 ( .A(n503), .B(n308), .Y(n42) );
  NAND2BX1 U756 ( .AN(n310), .B(n311), .Y(n43) );
  XOR2X1 U757 ( .A(n300), .B(n40), .Y(SUM[5]) );
  NAND2X1 U758 ( .A(n358), .B(n299), .Y(n40) );
  CLKINVX1 U759 ( .A(n298), .Y(n358) );
  NAND2X1 U760 ( .A(n359), .B(n303), .Y(n41) );
  CLKINVX1 U761 ( .A(n302), .Y(n359) );
  NAND2BX1 U762 ( .AN(n315), .B(n316), .Y(n44) );
  NOR2X2 U763 ( .A(B[36]), .B(A[38]), .Y(n84) );
  NOR2X2 U764 ( .A(B[36]), .B(A[39]), .Y(n75) );
  NOR2X2 U765 ( .A(B[36]), .B(A[37]), .Y(n95) );
  NAND2X1 U766 ( .A(n517), .B(n47), .Y(n2) );
  NOR2X2 U767 ( .A(B[33]), .B(A[33]), .Y(n131) );
  NOR2X2 U768 ( .A(B[23]), .B(A[23]), .Y(n209) );
  NOR2X2 U769 ( .A(B[17]), .B(A[17]), .Y(n239) );
  NOR2X2 U770 ( .A(B[13]), .B(A[13]), .Y(n261) );
  NAND2X1 U771 ( .A(B[36]), .B(A[38]), .Y(n85) );
  NAND2X1 U772 ( .A(B[36]), .B(A[39]), .Y(n76) );
  NAND2X1 U773 ( .A(B[36]), .B(A[37]), .Y(n96) );
  NAND2X1 U774 ( .A(B[24]), .B(A[24]), .Y(n203) );
  NAND2X1 U775 ( .A(B[23]), .B(A[23]), .Y(n210) );
  NAND2X1 U776 ( .A(B[33]), .B(A[33]), .Y(n132) );
  NAND2X1 U777 ( .A(B[29]), .B(A[29]), .Y(n159) );
  NAND2X1 U778 ( .A(B[19]), .B(A[19]), .Y(n229) );
  CLKINVX1 U779 ( .A(n45), .Y(SUM[0]) );
endmodule


module CONV ( clk, reset, busy, ready, iaddr, idata, cwr, caddr_wr, cdata_wr, 
        crd, caddr_rd, cdata_rd, csel );
  output [11:0] iaddr;
  input [19:0] idata;
  output [11:0] caddr_wr;
  output [19:0] cdata_wr;
  output [11:0] caddr_rd;
  input [19:0] cdata_rd;
  output [2:0] csel;
  input clk, reset, ready;
  output busy, cwr, crd;
  wire   n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, N53, N55,
         N61, N71, N78, N85, N89, N90, N94, N98, N102, N109, N111, N114, N124,
         N128, N144, N145, N146, N147, N148, N149, N175, N176, N177, N178,
         N179, N180, N363, mulTemp_43, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470,
         N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, N496, N497, N815, N816, N817, N818, N819, N820,
         N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831,
         N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842,
         N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853,
         N854, N855, N856, N857, N858, n24, n26, n29, n30, n34, n39, n41, n43,
         n45, n47, n78, n79, n80, n82, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n210, n213, n218, n219, n220, n224, n225, n229, n238, n239, n244,
         n245, n246, n247, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n391, n392, n393, n394, n395, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n426, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, \add_112_S2/carry[5] , \add_112_S2/carry[4] ,
         \add_112_S2/carry[3] , \add_99/carry[5] , \add_99/carry[4] ,
         \add_99/carry[3] , \r356/carry[5] , \r356/carry[4] , \r356/carry[3] ,
         \r356/carry[2] , \r354/carry[5] , \r354/carry[4] , \r354/carry[3] ,
         \r354/carry[2] , n527, n528, n529, n530, n972, n534, n535, n576, n966,
         n578, n967, n580, n969, n582, n970, n584, n971, n592, n968, n596,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n952, n954,
         n956, n958, n960, n962, n964;
  wire   [43:0] convTemp;
  wire   [20:1] roundTemp;
  wire   [5:0] index_X;
  wire   [5:0] index_X_Before;
  wire   [5:0] index_X_After;
  wire   [5:0] index_Y;
  wire   [5:0] index_Y_Before;
  wire   [5:0] index_Y_After;
  wire   [2:0] next_State;
  wire   [19:0] idataTemp;
  wire   [38:0] mulTemp;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign csel[2] = 1'b0;

  NOR2BX4 U88 ( .AN(n104), .B(n870), .Y(n84) );
  DFFRX1 \convTemp_reg[43]  ( .D(n440), .CK(clk), .RN(n650), .Q(convTemp[43]), 
        .QN(n346) );
  DFFRX1 \convTemp_reg[7]  ( .D(n476), .CK(clk), .RN(n649), .Q(convTemp[7]), 
        .QN(n310) );
  DFFRX1 \convTemp_reg[8]  ( .D(n475), .CK(clk), .RN(n649), .Q(convTemp[8]), 
        .QN(n311) );
  DFFRX1 \convTemp_reg[9]  ( .D(n474), .CK(clk), .RN(n649), .Q(convTemp[9]), 
        .QN(n312) );
  DFFRX1 \convTemp_reg[11]  ( .D(n472), .CK(clk), .RN(n649), .Q(convTemp[11]), 
        .QN(n314) );
  DFFRX1 \convTemp_reg[13]  ( .D(n470), .CK(clk), .RN(n648), .Q(convTemp[13]), 
        .QN(n316) );
  DFFRX2 \index_Y_reg[0]  ( .D(n520), .CK(clk), .RN(n654), .Q(N175), .QN(n402)
         );
  DFFRX1 \convTemp_reg[0]  ( .D(n483), .CK(clk), .RN(n650), .Q(convTemp[0]), 
        .QN(n303) );
  DFFRX1 \convTemp_reg[1]  ( .D(n482), .CK(clk), .RN(n649), .Q(convTemp[1]), 
        .QN(n304) );
  DFFRX1 \convTemp_reg[2]  ( .D(n481), .CK(clk), .RN(n649), .Q(convTemp[2]), 
        .QN(n305) );
  DFFRX1 \convTemp_reg[3]  ( .D(n480), .CK(clk), .RN(n649), .Q(convTemp[3]), 
        .QN(n306) );
  DFFRX1 \convTemp_reg[4]  ( .D(n479), .CK(clk), .RN(n649), .Q(convTemp[4]), 
        .QN(n307) );
  DFFRX1 \convTemp_reg[5]  ( .D(n478), .CK(clk), .RN(n649), .Q(convTemp[5]), 
        .QN(n308) );
  DFFRX1 \convTemp_reg[6]  ( .D(n477), .CK(clk), .RN(n649), .Q(convTemp[6]), 
        .QN(n309) );
  EDFFX1 \idataTemp_reg[16]  ( .D(idata[16]), .E(n529), .CK(clk), .Q(
        idataTemp[16]) );
  EDFFX1 \idataTemp_reg[10]  ( .D(idata[10]), .E(n529), .CK(clk), .Q(
        idataTemp[10]) );
  EDFFX1 \idataTemp_reg[8]  ( .D(idata[8]), .E(n529), .CK(clk), .Q(
        idataTemp[8]) );
  EDFFX1 \idataTemp_reg[6]  ( .D(idata[6]), .E(n529), .CK(clk), .Q(
        idataTemp[6]) );
  EDFFX1 \idataTemp_reg[4]  ( .D(idata[4]), .E(n529), .CK(clk), .Q(
        idataTemp[4]) );
  EDFFX1 \idataTemp_reg[2]  ( .D(idata[2]), .E(n529), .CK(clk), .Q(
        idataTemp[2]) );
  EDFFX1 \idataTemp_reg[17]  ( .D(idata[17]), .E(n529), .CK(clk), .Q(
        idataTemp[17]) );
  EDFFX1 \idataTemp_reg[13]  ( .D(idata[13]), .E(n529), .CK(clk), .Q(
        idataTemp[13]) );
  EDFFX1 \idataTemp_reg[11]  ( .D(idata[11]), .E(n529), .CK(clk), .Q(
        idataTemp[11]) );
  EDFFX1 \idataTemp_reg[9]  ( .D(idata[9]), .E(n529), .CK(clk), .Q(
        idataTemp[9]) );
  EDFFX1 \idataTemp_reg[7]  ( .D(idata[7]), .E(n529), .CK(clk), .Q(
        idataTemp[7]) );
  EDFFX1 \idataTemp_reg[5]  ( .D(idata[5]), .E(n529), .CK(clk), .Q(
        idataTemp[5]) );
  EDFFX1 \idataTemp_reg[0]  ( .D(idata[0]), .E(n529), .CK(clk), .Q(
        idataTemp[0]) );
  EDFFX1 \idataTemp_reg[15]  ( .D(idata[15]), .E(n529), .CK(clk), .Q(
        idataTemp[15]) );
  EDFFX1 \idataTemp_reg[1]  ( .D(idata[1]), .E(n529), .CK(clk), .Q(
        idataTemp[1]) );
  DFFRX1 \convTemp_reg[36]  ( .D(n447), .CK(clk), .RN(n647), .Q(convTemp[36]), 
        .QN(n339) );
  DFFRX1 \convTemp_reg[37]  ( .D(n446), .CK(clk), .RN(n647), .Q(convTemp[37]), 
        .QN(n340) );
  DFFRX1 \convTemp_reg[38]  ( .D(n445), .CK(clk), .RN(n646), .Q(convTemp[38]), 
        .QN(n341) );
  DFFRX1 \convTemp_reg[39]  ( .D(n444), .CK(clk), .RN(n646), .Q(convTemp[39]), 
        .QN(n342) );
  DFFRX1 \convTemp_reg[35]  ( .D(n448), .CK(clk), .RN(n650), .Q(convTemp[35]), 
        .QN(n338) );
  DFFRX1 \current_State_reg[0]  ( .D(next_State[0]), .CK(clk), .RN(n646), .Q(
        n866), .QN(n374) );
  DFFRX1 \index_Y_reg[3]  ( .D(n517), .CK(clk), .RN(n653), .Q(index_Y[3]), 
        .QN(n399) );
  DFFRX1 \index_X_reg[4]  ( .D(n511), .CK(clk), .RN(n654), .Q(index_X[4]), 
        .QN(n392) );
  DFFRX1 \index_X_reg[3]  ( .D(n512), .CK(clk), .RN(n654), .Q(index_X[3]), 
        .QN(n393) );
  DFFRX1 \index_X_reg[5]  ( .D(n521), .CK(clk), .RN(n654), .Q(index_X[5]), 
        .QN(n391) );
  DFFRX1 \index_Y_reg[5]  ( .D(n522), .CK(clk), .RN(n654), .Q(index_Y[5]), 
        .QN(n397) );
  DFFRX1 \index_Y_reg[4]  ( .D(n516), .CK(clk), .RN(n654), .Q(index_Y[4]), 
        .QN(n398) );
  DFFRX1 \index_X_reg[2]  ( .D(n513), .CK(clk), .RN(n654), .Q(index_X[2]), 
        .QN(n394) );
  DFFRX1 \index_X_reg[1]  ( .D(n514), .CK(clk), .RN(n654), .Q(index_X[1]), 
        .QN(n395) );
  DFFRX1 \convTemp_reg[19]  ( .D(n464), .CK(clk), .RN(n648), .Q(convTemp[19]), 
        .QN(n322) );
  DFFRX1 \convTemp_reg[31]  ( .D(n452), .CK(clk), .RN(n647), .Q(convTemp[31]), 
        .QN(n334) );
  DFFRX1 \convTemp_reg[33]  ( .D(n450), .CK(clk), .RN(n647), .Q(convTemp[33]), 
        .QN(n336) );
  DFFRX1 \index_Y_reg[1]  ( .D(n519), .CK(clk), .RN(n654), .Q(index_Y[1]), 
        .QN(n401) );
  DFFRX1 \index_Y_reg[2]  ( .D(n518), .CK(clk), .RN(n653), .Q(index_Y[2]), 
        .QN(n400) );
  DFFRX1 \convTemp_reg[15]  ( .D(n468), .CK(clk), .RN(n648), .Q(convTemp[15]), 
        .QN(n318) );
  DFFRX1 \convTemp_reg[17]  ( .D(n466), .CK(clk), .RN(n648), .Q(convTemp[17]), 
        .QN(n320) );
  DFFRX1 \convTemp_reg[26]  ( .D(n457), .CK(clk), .RN(n647), .Q(convTemp[26]), 
        .QN(n329) );
  DFFRX1 \convTemp_reg[29]  ( .D(n454), .CK(clk), .RN(n647), .Q(convTemp[29]), 
        .QN(n332) );
  DFFRX1 \convTemp_reg[25]  ( .D(n458), .CK(clk), .RN(n647), .Q(convTemp[25]), 
        .QN(n328) );
  DFFRX1 \convTemp_reg[28]  ( .D(n455), .CK(clk), .RN(n647), .Q(convTemp[28]), 
        .QN(n331) );
  DFFRX1 \convTemp_reg[21]  ( .D(n462), .CK(clk), .RN(n648), .Q(convTemp[21]), 
        .QN(n324) );
  DFFRX1 \convTemp_reg[23]  ( .D(n460), .CK(clk), .RN(n648), .Q(convTemp[23]), 
        .QN(n326) );
  DFFRX1 \convTemp_reg[24]  ( .D(n459), .CK(clk), .RN(n648), .Q(convTemp[24]), 
        .QN(n327) );
  DFFRX1 \current_State_reg[2]  ( .D(next_State[2]), .CK(clk), .RN(n646), .Q(
        n865), .QN(n423) );
  DFFRX4 \counterRead_reg[2]  ( .D(n523), .CK(clk), .RN(n646), .Q(n606), .QN(
        n426) );
  DFFRHQX8 \counterRead_reg[3]  ( .D(n525), .CK(clk), .RN(n646), .Q(n610) );
  DFFRX1 \convTemp_reg[14]  ( .D(n469), .CK(clk), .RN(n648), .Q(convTemp[14]), 
        .QN(n317) );
  DFFRX1 \convTemp_reg[12]  ( .D(n471), .CK(clk), .RN(n649), .Q(convTemp[12]), 
        .QN(n315) );
  DFFRX1 \convTemp_reg[34]  ( .D(n449), .CK(clk), .RN(n647), .Q(convTemp[34]), 
        .QN(n337) );
  DFFRX1 \convTemp_reg[10]  ( .D(n473), .CK(clk), .RN(n649), .Q(convTemp[10]), 
        .QN(n313) );
  DFFRX1 \convTemp_reg[30]  ( .D(n453), .CK(clk), .RN(n647), .Q(convTemp[30]), 
        .QN(n333) );
  DFFRX1 \convTemp_reg[18]  ( .D(n465), .CK(clk), .RN(n648), .Q(convTemp[18]), 
        .QN(n321) );
  DFFRX1 \convTemp_reg[22]  ( .D(n461), .CK(clk), .RN(n648), .Q(convTemp[22]), 
        .QN(n325) );
  DFFRX1 \convTemp_reg[16]  ( .D(n467), .CK(clk), .RN(n648), .Q(convTemp[16]), 
        .QN(n319) );
  DFFRX1 \convTemp_reg[40]  ( .D(n443), .CK(clk), .RN(n646), .Q(convTemp[40]), 
        .QN(n343) );
  DFFRX1 \convTemp_reg[41]  ( .D(n442), .CK(clk), .RN(n646), .Q(convTemp[41]), 
        .QN(n344) );
  DFFRX1 \convTemp_reg[42]  ( .D(n441), .CK(clk), .RN(n646), .Q(convTemp[42]), 
        .QN(n345) );
  DFFRX1 \convTemp_reg[27]  ( .D(n456), .CK(clk), .RN(n647), .Q(convTemp[27]), 
        .QN(n330) );
  DFFRHQX8 \counterRead_reg[1]  ( .D(n524), .CK(clk), .RN(n646), .Q(n608) );
  DFFRX2 \convTemp_reg[32]  ( .D(n451), .CK(clk), .RN(n647), .Q(convTemp[32]), 
        .QN(n335) );
  DFFRX1 \csel_reg[1]  ( .D(n508), .CK(clk), .RN(n653), .Q(n950), .QN(n596) );
  DFFRX1 crd_reg ( .D(n389), .CK(clk), .RN(n653), .Q(n937), .QN(n375) );
  DFFRX1 \caddr_wr_reg[0]  ( .D(n484), .CK(clk), .RN(n651), .Q(n916), .QN(n439) );
  DFFRX1 \caddr_wr_reg[1]  ( .D(n485), .CK(clk), .RN(n652), .Q(n915), .QN(n438) );
  DFFRX1 \caddr_wr_reg[2]  ( .D(n486), .CK(clk), .RN(n652), .Q(n914), .QN(n437) );
  DFFRX1 \caddr_wr_reg[3]  ( .D(n487), .CK(clk), .RN(n652), .Q(n913), .QN(n436) );
  DFFRX1 \caddr_wr_reg[4]  ( .D(n488), .CK(clk), .RN(n652), .Q(n912), .QN(n435) );
  DFFRX1 \caddr_wr_reg[5]  ( .D(n489), .CK(clk), .RN(n652), .Q(n911), .QN(n434) );
  DFFRX1 \caddr_wr_reg[6]  ( .D(n490), .CK(clk), .RN(n652), .Q(n910), .QN(n433) );
  DFFRX1 \caddr_wr_reg[7]  ( .D(n491), .CK(clk), .RN(n652), .Q(n909), .QN(n432) );
  DFFRX1 \caddr_wr_reg[8]  ( .D(n492), .CK(clk), .RN(n652), .Q(n908), .QN(n431) );
  DFFRX1 \caddr_wr_reg[9]  ( .D(n493), .CK(clk), .RN(n652), .Q(n907), .QN(n430) );
  DFFRX1 \caddr_rd_reg[0]  ( .D(n496), .CK(clk), .RN(n654), .Q(n949), .QN(n300) );
  DFFRX1 \caddr_rd_reg[1]  ( .D(n497), .CK(clk), .RN(n654), .Q(n948), .QN(n299) );
  DFFRX1 \caddr_rd_reg[2]  ( .D(n498), .CK(clk), .RN(n655), .Q(n947), .QN(n298) );
  DFFRX1 \caddr_rd_reg[3]  ( .D(n499), .CK(clk), .RN(n655), .Q(n946), .QN(n297) );
  DFFRX1 \caddr_rd_reg[4]  ( .D(n500), .CK(clk), .RN(n655), .Q(n945), .QN(n296) );
  DFFRX1 \caddr_rd_reg[5]  ( .D(n501), .CK(clk), .RN(n655), .Q(n944), .QN(n295) );
  DFFRX1 \caddr_rd_reg[6]  ( .D(n502), .CK(clk), .RN(n655), .Q(n943), .QN(n294) );
  DFFRX1 \caddr_rd_reg[7]  ( .D(n503), .CK(clk), .RN(n655), .Q(n942), .QN(n293) );
  DFFRX1 \caddr_rd_reg[8]  ( .D(n504), .CK(clk), .RN(n655), .Q(n941), .QN(n292) );
  DFFRX1 \caddr_rd_reg[9]  ( .D(n505), .CK(clk), .RN(n655), .Q(n940), .QN(n291) );
  DFFRX1 \caddr_rd_reg[10]  ( .D(n506), .CK(clk), .RN(n655), .Q(n939), .QN(
        n290) );
  DFFRX1 \caddr_rd_reg[11]  ( .D(n507), .CK(clk), .RN(n655), .Q(n938), .QN(
        n289) );
  DFFRX1 \csel_reg[0]  ( .D(n388), .CK(clk), .RN(n653), .Q(n951), .QN(n373) );
  DFFRX1 \caddr_wr_reg[10]  ( .D(n494), .CK(clk), .RN(n652), .Q(n906), .QN(
        n302) );
  DFFRX1 \caddr_wr_reg[11]  ( .D(n495), .CK(clk), .RN(n652), .Q(n905), .QN(
        n301) );
  DFFRX1 \iaddr_reg[0]  ( .D(n376), .CK(clk), .RN(n652), .Q(n904), .QN(n367)
         );
  DFFRX1 \iaddr_reg[1]  ( .D(n377), .CK(clk), .RN(n653), .Q(n903), .QN(n368)
         );
  DFFRX1 \iaddr_reg[2]  ( .D(n378), .CK(clk), .RN(n653), .Q(n902), .QN(n369)
         );
  DFFRX1 \iaddr_reg[3]  ( .D(n379), .CK(clk), .RN(n653), .Q(n901), .QN(n370)
         );
  DFFRX1 \iaddr_reg[4]  ( .D(n380), .CK(clk), .RN(n653), .Q(n900), .QN(n371)
         );
  DFFRX1 \iaddr_reg[5]  ( .D(n381), .CK(clk), .RN(n653), .Q(n899), .QN(n372)
         );
  DFFRX1 busy_reg ( .D(n510), .CK(clk), .RN(n653), .Q(n898), .QN(n429) );
  DFFRX1 \current_State_reg[1]  ( .D(next_State[1]), .CK(clk), .RN(n868), .Q(
        n660), .QN(n424) );
  EDFFXL \idataTemp_reg[19]  ( .D(idata[19]), .E(n529), .CK(clk), .Q(
        idataTemp[19]) );
  EDFFXL \idataTemp_reg[12]  ( .D(idata[12]), .E(n529), .CK(clk), .Q(
        idataTemp[12]) );
  EDFFXL \idataTemp_reg[18]  ( .D(idata[18]), .E(n529), .CK(clk), .Q(
        idataTemp[18]) );
  EDFFXL \idataTemp_reg[14]  ( .D(idata[14]), .E(n529), .CK(clk), .Q(
        idataTemp[14]) );
  DFFRX1 \convTemp_reg[20]  ( .D(n463), .CK(clk), .RN(n648), .Q(convTemp[20]), 
        .QN(n323) );
  DFFRHQX4 \counterRead_reg[0]  ( .D(n526), .CK(clk), .RN(n646), .Q(n603) );
  DFFRX1 \cdata_wr_reg[12]  ( .D(n415), .CK(clk), .RN(n651), .Q(n924), .QN(
        n359) );
  DFFRX1 \cdata_wr_reg[19]  ( .D(n422), .CK(clk), .RN(n651), .Q(n917), .QN(
        n366) );
  DFFRX1 \cdata_wr_reg[5]  ( .D(n408), .CK(clk), .RN(n650), .Q(n931), .QN(n352) );
  DFFRX1 \cdata_wr_reg[8]  ( .D(n411), .CK(clk), .RN(n650), .Q(n928), .QN(n355) );
  DFFRX1 \cdata_wr_reg[3]  ( .D(n406), .CK(clk), .RN(n650), .Q(n933), .QN(n350) );
  DFFRX1 \cdata_wr_reg[0]  ( .D(n403), .CK(clk), .RN(n651), .Q(n936), .QN(n347) );
  DFFRX1 \cdata_wr_reg[18]  ( .D(n421), .CK(clk), .RN(n651), .Q(n918), .QN(
        n365) );
  DFFRX1 \cdata_wr_reg[9]  ( .D(n412), .CK(clk), .RN(n650), .Q(n927), .QN(n356) );
  DFFRX1 \cdata_wr_reg[11]  ( .D(n414), .CK(clk), .RN(n651), .Q(n925), .QN(
        n358) );
  DFFRX1 \cdata_wr_reg[13]  ( .D(n416), .CK(clk), .RN(n651), .Q(n923), .QN(
        n360) );
  DFFRX1 \cdata_wr_reg[4]  ( .D(n407), .CK(clk), .RN(n650), .Q(n932), .QN(n351) );
  DFFRX1 \cdata_wr_reg[15]  ( .D(n418), .CK(clk), .RN(n651), .Q(n921), .QN(
        n362) );
  DFFRX1 \cdata_wr_reg[6]  ( .D(n409), .CK(clk), .RN(n650), .Q(n930), .QN(n353) );
  DFFRX1 \cdata_wr_reg[17]  ( .D(n420), .CK(clk), .RN(n651), .Q(n919), .QN(
        n364) );
  DFFRX1 \cdata_wr_reg[14]  ( .D(n417), .CK(clk), .RN(n651), .Q(n922), .QN(
        n361) );
  DFFRX1 \cdata_wr_reg[10]  ( .D(n413), .CK(clk), .RN(n651), .Q(n926), .QN(
        n357) );
  DFFRX1 \cdata_wr_reg[2]  ( .D(n405), .CK(clk), .RN(n650), .Q(n934), .QN(n349) );
  DFFRX1 \cdata_wr_reg[1]  ( .D(n404), .CK(clk), .RN(n650), .Q(n935), .QN(n348) );
  DFFRX1 \cdata_wr_reg[7]  ( .D(n410), .CK(clk), .RN(n650), .Q(n929), .QN(n354) );
  DFFRX1 \cdata_wr_reg[16]  ( .D(n419), .CK(clk), .RN(n651), .Q(n920), .QN(
        n363) );
  EDFFX2 \idataTemp_reg[3]  ( .D(idata[3]), .E(n529), .CK(clk), .Q(
        idataTemp[3]) );
  INVX4 U421 ( .A(n839), .Y(n850) );
  BUFX4 U422 ( .A(mulTemp[6]), .Y(n527) );
  INVX3 U423 ( .A(n680), .Y(n672) );
  NAND2X2 U424 ( .A(n605), .B(n675), .Y(n837) );
  NAND2X1 U425 ( .A(n687), .B(n603), .Y(n673) );
  INVX3 U426 ( .A(n616), .Y(n630) );
  INVX8 U427 ( .A(n603), .Y(n604) );
  CLKAND2X6 U428 ( .A(n609), .B(n603), .Y(n605) );
  NAND2X6 U429 ( .A(n604), .B(n608), .Y(n674) );
  NAND2X1 U430 ( .A(n528), .B(n609), .Y(n683) );
  NAND2BX2 U431 ( .AN(n674), .B(n607), .Y(n681) );
  CLKINVX1 U432 ( .A(n707), .Y(n693) );
  NAND2X2 U433 ( .A(n676), .B(n849), .Y(n839) );
  AND2X2 U434 ( .A(n694), .B(n853), .Y(n614) );
  NAND2X4 U435 ( .A(n604), .B(n528), .Y(n707) );
  CLKBUFX3 U436 ( .A(n631), .Y(n632) );
  NOR2BX1 U437 ( .AN(n104), .B(n870), .Y(n631) );
  INVX3 U438 ( .A(n617), .Y(n629) );
  OAI2BB2XL U439 ( .B0(n870), .B1(n104), .A0N(n869), .A1N(n870), .Y(n617) );
  INVX3 U440 ( .A(n606), .Y(n607) );
  BUFX4 U441 ( .A(mulTemp[15]), .Y(n534) );
  CLKINVX1 U442 ( .A(n832), .Y(n717) );
  OAI31XL U443 ( .A0(n702), .A1(n701), .A2(n700), .B0(n624), .Y(n830) );
  OAI21XL U444 ( .A0(n363), .A1(n629), .B0(n100), .Y(n419) );
  AOI22X1 U445 ( .A0(roundTemp[17]), .A1(n626), .B0(cdata_rd[16]), .B1(n632), 
        .Y(n100) );
  OAI21XL U446 ( .A0(n354), .A1(n630), .B0(n91), .Y(n410) );
  AOI22X1 U447 ( .A0(roundTemp[8]), .A1(n625), .B0(cdata_rd[7]), .B1(n633), 
        .Y(n91) );
  OAI21XL U448 ( .A0(n348), .A1(n630), .B0(n85), .Y(n404) );
  AOI22X1 U449 ( .A0(roundTemp[2]), .A1(n625), .B0(cdata_rd[1]), .B1(n633), 
        .Y(n85) );
  OAI21XL U450 ( .A0(n349), .A1(n629), .B0(n86), .Y(n405) );
  AOI22X1 U451 ( .A0(roundTemp[3]), .A1(n625), .B0(cdata_rd[2]), .B1(n632), 
        .Y(n86) );
  OAI21XL U452 ( .A0(n357), .A1(n629), .B0(n94), .Y(n413) );
  AOI22X1 U453 ( .A0(roundTemp[11]), .A1(n626), .B0(cdata_rd[10]), .B1(n632), 
        .Y(n94) );
  OAI21XL U454 ( .A0(n361), .A1(n629), .B0(n98), .Y(n417) );
  AOI22X1 U455 ( .A0(roundTemp[15]), .A1(n626), .B0(cdata_rd[14]), .B1(n632), 
        .Y(n98) );
  OAI21XL U456 ( .A0(n364), .A1(n630), .B0(n101), .Y(n420) );
  AOI22X1 U457 ( .A0(roundTemp[18]), .A1(n626), .B0(cdata_rd[17]), .B1(n633), 
        .Y(n101) );
  OAI21XL U458 ( .A0(n353), .A1(n629), .B0(n90), .Y(n409) );
  AOI22X1 U459 ( .A0(roundTemp[7]), .A1(n625), .B0(cdata_rd[6]), .B1(n632), 
        .Y(n90) );
  OAI21XL U460 ( .A0(n362), .A1(n630), .B0(n99), .Y(n418) );
  AOI22X1 U461 ( .A0(roundTemp[16]), .A1(n626), .B0(cdata_rd[15]), .B1(n633), 
        .Y(n99) );
  OAI21XL U462 ( .A0(n351), .A1(n629), .B0(n88), .Y(n407) );
  AOI22X1 U463 ( .A0(roundTemp[5]), .A1(n625), .B0(cdata_rd[4]), .B1(n632), 
        .Y(n88) );
  OAI21XL U464 ( .A0(n360), .A1(n630), .B0(n97), .Y(n416) );
  AOI22X1 U465 ( .A0(roundTemp[14]), .A1(n626), .B0(cdata_rd[13]), .B1(n633), 
        .Y(n97) );
  OAI21XL U466 ( .A0(n358), .A1(n630), .B0(n95), .Y(n414) );
  AOI22X1 U467 ( .A0(roundTemp[12]), .A1(n626), .B0(cdata_rd[11]), .B1(n633), 
        .Y(n95) );
  OAI21XL U468 ( .A0(n356), .A1(n630), .B0(n93), .Y(n412) );
  AOI22X1 U469 ( .A0(roundTemp[10]), .A1(n625), .B0(cdata_rd[9]), .B1(n633), 
        .Y(n93) );
  OAI21XL U470 ( .A0(n365), .A1(n629), .B0(n102), .Y(n421) );
  AOI22X1 U471 ( .A0(roundTemp[19]), .A1(n626), .B0(cdata_rd[18]), .B1(n632), 
        .Y(n102) );
  OAI21XL U472 ( .A0(n347), .A1(n629), .B0(n82), .Y(n403) );
  AOI22X1 U473 ( .A0(roundTemp[1]), .A1(n625), .B0(cdata_rd[0]), .B1(n632), 
        .Y(n82) );
  OAI21XL U474 ( .A0(n350), .A1(n630), .B0(n87), .Y(n406) );
  AOI22X1 U475 ( .A0(roundTemp[4]), .A1(n625), .B0(cdata_rd[3]), .B1(n633), 
        .Y(n87) );
  OAI21XL U476 ( .A0(n355), .A1(n629), .B0(n92), .Y(n411) );
  AOI22X1 U477 ( .A0(roundTemp[9]), .A1(n625), .B0(cdata_rd[8]), .B1(n632), 
        .Y(n92) );
  OAI21XL U478 ( .A0(n352), .A1(n630), .B0(n89), .Y(n408) );
  AOI22X1 U479 ( .A0(roundTemp[6]), .A1(n625), .B0(cdata_rd[5]), .B1(n633), 
        .Y(n89) );
  OAI21XL U480 ( .A0(n366), .A1(n630), .B0(n103), .Y(n422) );
  AOI22X1 U481 ( .A0(roundTemp[20]), .A1(n626), .B0(cdata_rd[19]), .B1(n633), 
        .Y(n103) );
  OAI21XL U482 ( .A0(n359), .A1(n629), .B0(n96), .Y(n415) );
  AOI22X1 U483 ( .A0(roundTemp[13]), .A1(n626), .B0(cdata_rd[12]), .B1(n632), 
        .Y(n96) );
  CLKINVX1 U484 ( .A(n605), .Y(n670) );
  AND2X6 U485 ( .A(n426), .B(n610), .Y(n528) );
  INVXL U486 ( .A(mulTemp[36]), .Y(n722) );
  CLKAND2X3 U487 ( .A(n624), .B(n656), .Y(n529) );
  AND2X2 U488 ( .A(n639), .B(n708), .Y(n530) );
  CLKINVX1 U489 ( .A(n848), .Y(n676) );
  OAI211X4 U492 ( .A0(n604), .A1(n851), .B0(n683), .C0(n682), .Y(N114) );
  INVX6 U493 ( .A(n608), .Y(n609) );
  INVX6 U494 ( .A(n851), .Y(n675) );
  OR2X2 U495 ( .A(n610), .B(n426), .Y(n851) );
  BUFX6 U496 ( .A(n611), .Y(n535) );
  INVXL U497 ( .A(n610), .Y(n611) );
  NAND2X4 U498 ( .A(n675), .B(n608), .Y(n853) );
  NAND3BXL U499 ( .AN(n693), .B(n618), .C(n681), .Y(N78) );
  INVX8 U500 ( .A(n681), .Y(N55) );
  NAND2X1 U501 ( .A(n849), .B(n608), .Y(n682) );
  BUFX12 U502 ( .A(n920), .Y(cdata_wr[16]) );
  BUFX12 U503 ( .A(n929), .Y(cdata_wr[7]) );
  BUFX12 U504 ( .A(n935), .Y(cdata_wr[1]) );
  BUFX12 U505 ( .A(n934), .Y(cdata_wr[2]) );
  BUFX12 U506 ( .A(n926), .Y(cdata_wr[10]) );
  BUFX12 U507 ( .A(n922), .Y(cdata_wr[14]) );
  BUFX12 U508 ( .A(n919), .Y(cdata_wr[17]) );
  BUFX12 U509 ( .A(n898), .Y(busy) );
  BUFX12 U510 ( .A(n899), .Y(iaddr[5]) );
  BUFX12 U511 ( .A(n900), .Y(iaddr[4]) );
  BUFX12 U512 ( .A(n901), .Y(iaddr[3]) );
  BUFX12 U513 ( .A(n902), .Y(iaddr[2]) );
  BUFX12 U514 ( .A(n903), .Y(iaddr[1]) );
  BUFX12 U515 ( .A(n904), .Y(iaddr[0]) );
  BUFX12 U516 ( .A(n905), .Y(caddr_wr[11]) );
  BUFX12 U517 ( .A(n906), .Y(caddr_wr[10]) );
  BUFX12 U518 ( .A(n951), .Y(csel[0]) );
  BUFX12 U519 ( .A(n938), .Y(caddr_rd[11]) );
  BUFX12 U520 ( .A(n939), .Y(caddr_rd[10]) );
  BUFX12 U521 ( .A(n940), .Y(caddr_rd[9]) );
  BUFX12 U522 ( .A(n941), .Y(caddr_rd[8]) );
  BUFX12 U523 ( .A(n942), .Y(caddr_rd[7]) );
  BUFX12 U524 ( .A(n943), .Y(caddr_rd[6]) );
  BUFX12 U525 ( .A(n944), .Y(caddr_rd[5]) );
  BUFX12 U526 ( .A(n945), .Y(caddr_rd[4]) );
  BUFX12 U527 ( .A(n946), .Y(caddr_rd[3]) );
  BUFX12 U528 ( .A(n947), .Y(caddr_rd[2]) );
  BUFX12 U529 ( .A(n948), .Y(caddr_rd[1]) );
  BUFX12 U530 ( .A(n949), .Y(caddr_rd[0]) );
  BUFX12 U531 ( .A(n907), .Y(caddr_wr[9]) );
  BUFX12 U532 ( .A(n908), .Y(caddr_wr[8]) );
  BUFX12 U533 ( .A(n909), .Y(caddr_wr[7]) );
  BUFX12 U534 ( .A(n910), .Y(caddr_wr[6]) );
  BUFX12 U535 ( .A(n911), .Y(caddr_wr[5]) );
  BUFX12 U536 ( .A(n912), .Y(caddr_wr[4]) );
  BUFX12 U537 ( .A(n913), .Y(caddr_wr[3]) );
  BUFX12 U538 ( .A(n914), .Y(caddr_wr[2]) );
  BUFX12 U539 ( .A(n915), .Y(caddr_wr[1]) );
  BUFX12 U540 ( .A(n916), .Y(caddr_wr[0]) );
  BUFX12 U541 ( .A(n937), .Y(crd) );
  BUFX12 U547 ( .A(n930), .Y(cdata_wr[6]) );
  BUFX12 U548 ( .A(n921), .Y(cdata_wr[15]) );
  BUFX12 U549 ( .A(n932), .Y(cdata_wr[4]) );
  BUFX12 U550 ( .A(n923), .Y(cdata_wr[13]) );
  BUFX12 U551 ( .A(n925), .Y(cdata_wr[11]) );
  BUFX12 U552 ( .A(n927), .Y(cdata_wr[9]) );
  BUFX12 U554 ( .A(n918), .Y(cdata_wr[18]) );
  BUFX12 U555 ( .A(n936), .Y(cdata_wr[0]) );
  INVX12 U556 ( .A(n596), .Y(csel[1]) );
  BUFX12 U557 ( .A(n933), .Y(cdata_wr[3]) );
  BUFX12 U558 ( .A(n928), .Y(cdata_wr[8]) );
  BUFX12 U559 ( .A(n931), .Y(cdata_wr[5]) );
  BUFX12 U560 ( .A(n917), .Y(cdata_wr[19]) );
  BUFX12 U561 ( .A(n924), .Y(cdata_wr[12]) );
  NAND2X2 U562 ( .A(n683), .B(n707), .Y(n680) );
  NAND3BXL U563 ( .AN(n850), .B(n707), .C(n684), .Y(N128) );
  INVXL U564 ( .A(mulTemp[31]), .Y(n734) );
  NAND2X4 U565 ( .A(n603), .B(n608), .Y(n848) );
  CLKINVX8 U566 ( .A(n688), .Y(n849) );
  NAND2X6 U567 ( .A(n535), .B(n607), .Y(n688) );
  INVXL U568 ( .A(mulTemp[21]), .Y(n764) );
  NAND2X1 U569 ( .A(n684), .B(n678), .Y(N102) );
  BUFX20 U570 ( .A(n84), .Y(n633) );
  AOI2BB1XL U571 ( .A0N(n688), .A1N(n608), .B0(n687), .Y(n689) );
  INVX3 U572 ( .A(n853), .Y(n687) );
  NAND2X2 U573 ( .A(n882), .B(n609), .Y(n705) );
  NAND2X8 U574 ( .A(n604), .B(n675), .Y(n684) );
  NAND3X1 U575 ( .A(n612), .B(n832), .C(n831), .Y(n440) );
  AOI22X1 U576 ( .A0(N497), .A1(n530), .B0(N858), .B1(n613), .Y(n612) );
  OR2XL U577 ( .A(n689), .B(n603), .Y(n840) );
  NAND2X6 U578 ( .A(n605), .B(n528), .Y(n694) );
  OAI2BB1XL U579 ( .A0N(n676), .A1N(n535), .B0(n854), .Y(n677) );
  NAND2X2 U580 ( .A(n693), .B(n609), .Y(n854) );
  INVXL U581 ( .A(mulTemp[35]), .Y(n833) );
  INVXL U582 ( .A(mulTemp[27]), .Y(n746) );
  NAND2XL U583 ( .A(n618), .B(n694), .Y(N71) );
  NAND2X4 U584 ( .A(n705), .B(n619), .Y(N124) );
  AO21XL U585 ( .A0(n687), .A1(n604), .B0(n679), .Y(N109) );
  INVXL U586 ( .A(n694), .Y(n679) );
  AO21XL U587 ( .A0(n535), .A1(n608), .B0(n680), .Y(N111) );
  INVX1 U588 ( .A(mulTemp[20]), .Y(n767) );
  INVXL U589 ( .A(mulTemp[33]), .Y(n728) );
  INVXL U590 ( .A(mulTemp[29]), .Y(n740) );
  INVX1 U591 ( .A(mulTemp[32]), .Y(n731) );
  INVX1 U592 ( .A(mulTemp[30]), .Y(n737) );
  INVX1 U593 ( .A(mulTemp[34]), .Y(n725) );
  INVXL U594 ( .A(mulTemp[26]), .Y(n749) );
  INVXL U595 ( .A(mulTemp[25]), .Y(n752) );
  INVXL U596 ( .A(mulTemp[24]), .Y(n755) );
  INVXL U597 ( .A(mulTemp[28]), .Y(n743) );
  CLKINVX1 U598 ( .A(n830), .Y(n834) );
  INVX3 U599 ( .A(n266), .Y(n869) );
  NAND2XL U600 ( .A(n605), .B(n849), .Y(n838) );
  NAND3BX2 U601 ( .AN(n882), .B(n681), .C(n614), .Y(N89) );
  OAI2BB2X2 U602 ( .B0(n870), .B1(n104), .A0N(n869), .A1N(n870), .Y(n616) );
  NAND4XL U603 ( .A(n707), .B(n706), .C(n705), .D(n614), .Y(n708) );
  INVXL U604 ( .A(N85), .Y(n706) );
  OAI211XL U605 ( .A0(n696), .A1(n854), .B0(n695), .C0(n694), .Y(n698) );
  NAND3BXL U606 ( .AN(n883), .B(n693), .C(n608), .Y(n695) );
  NAND2X1 U607 ( .A(n268), .B(N144), .Y(n218) );
  AO22XL U608 ( .A0(n665), .A1(n699), .B0(n664), .B1(n610), .Y(n525) );
  NOR2X1 U609 ( .A(n866), .B(n79), .Y(n266) );
  NAND3BXL U610 ( .AN(n622), .B(n849), .C(n848), .Y(n856) );
  AND2X1 U611 ( .A(n849), .B(n627), .Y(n620) );
  AOI2BB1XL U612 ( .A0N(n851), .A1N(n608), .B0(n850), .Y(n852) );
  NAND2XL U613 ( .A(N55), .B(n535), .Y(n685) );
  INVXL U614 ( .A(mulTemp[19]), .Y(n770) );
  INVXL U615 ( .A(mulTemp[17]), .Y(n776) );
  INVXL U616 ( .A(mulTemp[18]), .Y(n773) );
  INVXL U617 ( .A(mulTemp[16]), .Y(n779) );
  INVXL U618 ( .A(n534), .Y(n782) );
  INVXL U619 ( .A(mulTemp[13]), .Y(n788) );
  INVXL U620 ( .A(mulTemp[14]), .Y(n785) );
  INVXL U621 ( .A(mulTemp[12]), .Y(n791) );
  INVXL U622 ( .A(mulTemp[9]), .Y(n800) );
  INVXL U623 ( .A(mulTemp[11]), .Y(n794) );
  INVXL U624 ( .A(mulTemp[10]), .Y(n797) );
  INVXL U625 ( .A(mulTemp[8]), .Y(n803) );
  INVXL U626 ( .A(mulTemp[7]), .Y(n806) );
  INVXL U627 ( .A(n527), .Y(n809) );
  INVXL U628 ( .A(mulTemp[5]), .Y(n812) );
  INVXL U629 ( .A(mulTemp[4]), .Y(n815) );
  INVXL U630 ( .A(mulTemp[3]), .Y(n818) );
  AOI2BB1XL U631 ( .A0N(n424), .A1N(n705), .B0(n704), .Y(n662) );
  CLKBUFX3 U632 ( .A(n229), .Y(n627) );
  MX2XL U633 ( .A(n666), .B(n665), .S0(n604), .Y(n526) );
  MX2XL U634 ( .A(n664), .B(n663), .S0(n607), .Y(n523) );
  AND2XL U635 ( .A(n665), .B(n676), .Y(n663) );
  NAND3X1 U636 ( .A(n865), .B(n866), .C(n424), .Y(n29) );
  ADDHXL U637 ( .A(index_Y[1]), .B(N175), .CO(\r356/carry[2] ), .S(
        index_Y_After[1]) );
  ADDHXL U638 ( .A(index_X[1]), .B(N144), .CO(\r354/carry[2] ), .S(
        index_X_After[1]) );
  ADDHXL U639 ( .A(index_Y[2]), .B(\r356/carry[2] ), .CO(\r356/carry[3] ), .S(
        index_Y_After[2]) );
  ADDHXL U640 ( .A(index_X[2]), .B(\r354/carry[2] ), .CO(\r354/carry[3] ), .S(
        index_X_After[2]) );
  ADDHXL U641 ( .A(index_Y[3]), .B(\r356/carry[3] ), .CO(\r356/carry[4] ), .S(
        index_Y_After[3]) );
  ADDHXL U642 ( .A(index_X[3]), .B(\r354/carry[3] ), .CO(\r354/carry[4] ), .S(
        index_X_After[3]) );
  ADDHXL U643 ( .A(index_Y[4]), .B(\r356/carry[4] ), .CO(\r356/carry[5] ), .S(
        index_Y_After[4]) );
  ADDHXL U644 ( .A(index_X[4]), .B(\r354/carry[4] ), .CO(\r354/carry[5] ), .S(
        index_X_After[4]) );
  CLKINVX1 U645 ( .A(mulTemp[23]), .Y(n758) );
  CLKINVX1 U646 ( .A(mulTemp[22]), .Y(n761) );
  NAND2X1 U647 ( .A(mulTemp_43), .B(n615), .Y(n832) );
  CLKBUFX3 U648 ( .A(n613), .Y(n638) );
  CLKBUFX3 U649 ( .A(n613), .Y(n637) );
  CLKINVX1 U650 ( .A(mulTemp[2]), .Y(n821) );
  NAND2X1 U651 ( .A(n837), .B(n839), .Y(N85) );
  AND2X2 U652 ( .A(n704), .B(n639), .Y(n613) );
  CLKBUFX3 U653 ( .A(n834), .Y(n639) );
  INVX3 U654 ( .A(n615), .Y(n634) );
  INVX3 U655 ( .A(n615), .Y(n635) );
  INVX3 U656 ( .A(n615), .Y(n636) );
  CLKINVX1 U657 ( .A(n837), .Y(n692) );
  CLKBUFX3 U658 ( .A(n834), .Y(n640) );
  CLKINVX1 U659 ( .A(mulTemp[1]), .Y(n824) );
  CLKINVX1 U660 ( .A(mulTemp[0]), .Y(n827) );
  CLKBUFX3 U661 ( .A(n645), .Y(n647) );
  CLKBUFX3 U662 ( .A(n645), .Y(n648) );
  CLKBUFX3 U663 ( .A(n645), .Y(n649) );
  CLKBUFX3 U664 ( .A(n645), .Y(n650) );
  CLKBUFX3 U665 ( .A(n645), .Y(n651) );
  CLKBUFX3 U666 ( .A(n645), .Y(n652) );
  CLKBUFX3 U667 ( .A(n645), .Y(n655) );
  CLKBUFX3 U668 ( .A(n645), .Y(n653) );
  CLKBUFX3 U669 ( .A(n645), .Y(n654) );
  CLKBUFX3 U670 ( .A(n645), .Y(n646) );
  NAND2X1 U671 ( .A(n853), .B(n672), .Y(N53) );
  CLKBUFX3 U672 ( .A(n509), .Y(n628) );
  NAND2X1 U673 ( .A(n869), .B(n623), .Y(n509) );
  CLKBUFX3 U674 ( .A(n643), .Y(n656) );
  CLKBUFX3 U675 ( .A(n644), .Y(n643) );
  AND2X2 U676 ( .A(n639), .B(n703), .Y(n615) );
  CLKINVX1 U677 ( .A(n673), .Y(n699) );
  CLKBUFX3 U678 ( .A(n530), .Y(n642) );
  CLKBUFX3 U679 ( .A(n530), .Y(n641) );
  NOR2BX2 U680 ( .AN(n257), .B(n869), .Y(n260) );
  NAND2X1 U681 ( .A(n618), .B(n838), .Y(n842) );
  CLKINVX1 U682 ( .A(n690), .Y(n704) );
  CLKINVX1 U683 ( .A(n667), .Y(n666) );
  CLKINVX1 U684 ( .A(n218), .Y(n883) );
  AO21X1 U685 ( .A0(n665), .A1(n848), .B0(n666), .Y(n664) );
  NAND2X1 U686 ( .A(n619), .B(n837), .Y(n843) );
  NAND2X1 U687 ( .A(n840), .B(n839), .Y(n841) );
  CLKINVX1 U688 ( .A(n856), .Y(n862) );
  NAND2X1 U689 ( .A(n266), .B(n218), .Y(n249) );
  NAND2X1 U690 ( .A(n853), .B(n678), .Y(N94) );
  CLKINVX1 U691 ( .A(n684), .Y(n882) );
  AND2X2 U692 ( .A(n673), .B(n705), .Y(n618) );
  AND2X2 U693 ( .A(n685), .B(n854), .Y(n619) );
  OAI211X1 U694 ( .A0(n610), .A1(n674), .B0(n672), .C0(n682), .Y(N61) );
  NAND3BX1 U695 ( .AN(n693), .B(n684), .C(n853), .Y(N90) );
  NAND2X1 U696 ( .A(n854), .B(n682), .Y(N98) );
  CLKBUFX3 U697 ( .A(n225), .Y(n623) );
  NAND2X1 U698 ( .A(next_State[2]), .B(next_State[0]), .Y(n225) );
  CLKBUFX3 U699 ( .A(n868), .Y(n644) );
  AND2X2 U700 ( .A(n692), .B(n210), .Y(n701) );
  AO22X1 U701 ( .A0(n699), .A1(n218), .B0(n698), .B1(n697), .Y(n700) );
  OAI211X1 U702 ( .A0(n213), .A1(n691), .B0(n690), .C0(n840), .Y(n702) );
  AOI221XL U703 ( .A0(n686), .A1(n218), .B0(n210), .B1(n703), .C0(n850), .Y(
        n691) );
  CLKINVX1 U704 ( .A(n210), .Y(n696) );
  CLKINVX1 U705 ( .A(n705), .Y(n686) );
  CLKINVX1 U706 ( .A(n685), .Y(n703) );
  OAI22X2 U707 ( .A0(n245), .A1(n29), .B0(n218), .B1(n869), .Y(n257) );
  NOR2BX2 U708 ( .AN(n257), .B(n29), .Y(n259) );
  NAND2X1 U709 ( .A(n528), .B(n676), .Y(n690) );
  NAND3BX1 U710 ( .AN(n627), .B(n690), .C(n668), .Y(n667) );
  CLKINVX1 U711 ( .A(n668), .Y(n665) );
  AO22X1 U712 ( .A0(n80), .A1(n865), .B0(n686), .B1(n627), .Y(next_State[2])
         );
  CLKBUFX3 U713 ( .A(n867), .Y(n624) );
  CLKINVX1 U714 ( .A(n622), .Y(n867) );
  CLKINVX1 U715 ( .A(n30), .Y(n697) );
  NAND2X1 U716 ( .A(n620), .B(n603), .Y(n844) );
  NAND2X1 U717 ( .A(n620), .B(n608), .Y(n846) );
  NOR2BX2 U718 ( .AN(n245), .B(n29), .Y(n252) );
  INVX3 U719 ( .A(n627), .Y(n870) );
  NAND2X1 U720 ( .A(n29), .B(n869), .Y(n250) );
  AO21X1 U721 ( .A0(n854), .A1(n853), .B0(n622), .Y(n864) );
  OR2X1 U722 ( .A(n622), .B(n852), .Y(n861) );
  CLKINVX1 U723 ( .A(index_Y_After[5]), .Y(n892) );
  CLKINVX1 U724 ( .A(index_X_After[5]), .Y(n884) );
  CLKBUFX3 U725 ( .A(n621), .Y(n626) );
  CLKBUFX3 U726 ( .A(n621), .Y(n625) );
  CLKINVX1 U727 ( .A(index_Y_After[1]), .Y(n897) );
  CLKINVX1 U728 ( .A(index_X_After[1]), .Y(n888) );
  CLKINVX1 U729 ( .A(index_Y_After[4]), .Y(n894) );
  CLKINVX1 U730 ( .A(index_Y_After[2]), .Y(n896) );
  CLKINVX1 U731 ( .A(index_Y_After[3]), .Y(n895) );
  CLKINVX1 U732 ( .A(index_X_After[4]), .Y(n885) );
  CLKINVX1 U733 ( .A(index_X_After[2]), .Y(n887) );
  CLKINVX1 U734 ( .A(index_X_After[3]), .Y(n886) );
  CLKBUFX3 U735 ( .A(n868), .Y(n645) );
  CLKINVX1 U736 ( .A(n838), .Y(n671) );
  NAND3BX1 U737 ( .AN(n717), .B(n714), .C(n713), .Y(n443) );
  NAND2X1 U738 ( .A(N855), .B(n613), .Y(n714) );
  AOI2BB2X1 U739 ( .B0(N494), .B1(n641), .A0N(n343), .A1N(n640), .Y(n713) );
  NAND2X1 U740 ( .A(n830), .B(convTemp[43]), .Y(n831) );
  NAND3BX1 U741 ( .AN(n717), .B(n710), .C(n709), .Y(n441) );
  NAND2X1 U742 ( .A(N857), .B(n613), .Y(n710) );
  AOI2BB2X1 U743 ( .B0(N496), .B1(n530), .A0N(n345), .A1N(n639), .Y(n709) );
  NAND3BX1 U744 ( .AN(n717), .B(n712), .C(n711), .Y(n442) );
  NAND2X1 U745 ( .A(N856), .B(n613), .Y(n712) );
  AOI2BB2X1 U746 ( .B0(N495), .B1(n642), .A0N(n344), .A1N(n640), .Y(n711) );
  CLKINVX1 U747 ( .A(n677), .Y(n678) );
  NAND3BX1 U748 ( .AN(n717), .B(n716), .C(n715), .Y(n444) );
  NAND2X1 U749 ( .A(N854), .B(n613), .Y(n716) );
  AOI2BB2X1 U750 ( .B0(N493), .B1(n641), .A0N(n342), .A1N(n640), .Y(n715) );
  NAND2X1 U751 ( .A(n727), .B(n726), .Y(n449) );
  AOI2BB2X1 U752 ( .B0(N849), .B1(n638), .A0N(n634), .A1N(n725), .Y(n727) );
  AOI2BB2X1 U753 ( .B0(N488), .B1(n642), .A0N(n337), .A1N(n834), .Y(n726) );
  NAND2X1 U754 ( .A(n736), .B(n735), .Y(n452) );
  AOI2BB2X1 U755 ( .B0(N846), .B1(n638), .A0N(n634), .A1N(n734), .Y(n736) );
  AOI2BB2X1 U756 ( .B0(N485), .B1(n642), .A0N(n334), .A1N(n640), .Y(n735) );
  NAND2X1 U757 ( .A(n739), .B(n738), .Y(n453) );
  AOI2BB2X1 U758 ( .B0(N845), .B1(n638), .A0N(n634), .A1N(n737), .Y(n739) );
  AOI2BB2X1 U759 ( .B0(N484), .B1(n642), .A0N(n333), .A1N(n640), .Y(n738) );
  NAND2X1 U760 ( .A(n742), .B(n741), .Y(n454) );
  AOI2BB2X1 U761 ( .B0(N844), .B1(n638), .A0N(n634), .A1N(n740), .Y(n742) );
  AOI2BB2X1 U762 ( .B0(N483), .B1(n642), .A0N(n332), .A1N(n640), .Y(n741) );
  NAND2X1 U763 ( .A(n745), .B(n744), .Y(n455) );
  AOI2BB2X1 U764 ( .B0(N843), .B1(n638), .A0N(n634), .A1N(n743), .Y(n745) );
  AOI2BB2X1 U765 ( .B0(N482), .B1(n642), .A0N(n331), .A1N(n639), .Y(n744) );
  NAND2X1 U766 ( .A(n760), .B(n759), .Y(n460) );
  AOI2BB2X1 U767 ( .B0(N838), .B1(n638), .A0N(n635), .A1N(n758), .Y(n760) );
  AOI2BB2X1 U768 ( .B0(N477), .B1(n642), .A0N(n326), .A1N(n640), .Y(n759) );
  NAND2X1 U769 ( .A(n719), .B(n718), .Y(n445) );
  AOI2BB2X1 U770 ( .B0(N853), .B1(n613), .A0N(n634), .A1N(n722), .Y(n719) );
  AOI2BB2X1 U771 ( .B0(N492), .B1(n641), .A0N(n341), .A1N(n834), .Y(n718) );
  NAND2X1 U772 ( .A(n721), .B(n720), .Y(n446) );
  AOI2BB2X1 U773 ( .B0(N852), .B1(n613), .A0N(n634), .A1N(n722), .Y(n721) );
  AOI2BB2X1 U774 ( .B0(N491), .B1(n642), .A0N(n340), .A1N(n834), .Y(n720) );
  NAND2X1 U775 ( .A(n724), .B(n723), .Y(n447) );
  AOI2BB2X1 U776 ( .B0(N851), .B1(n613), .A0N(n634), .A1N(n722), .Y(n724) );
  AOI2BB2X1 U777 ( .B0(N490), .B1(n641), .A0N(n339), .A1N(n639), .Y(n723) );
  NAND2X1 U778 ( .A(n836), .B(n835), .Y(n448) );
  AOI2BB2X1 U779 ( .B0(N850), .B1(n637), .A0N(n634), .A1N(n833), .Y(n836) );
  AOI2BB2X1 U780 ( .B0(N489), .B1(n641), .A0N(n338), .A1N(n640), .Y(n835) );
  NAND2X1 U781 ( .A(n730), .B(n729), .Y(n450) );
  AOI2BB2X1 U782 ( .B0(N848), .B1(n638), .A0N(n634), .A1N(n728), .Y(n730) );
  AOI2BB2X1 U783 ( .B0(N487), .B1(n642), .A0N(n336), .A1N(n639), .Y(n729) );
  NAND2X1 U784 ( .A(n748), .B(n747), .Y(n456) );
  AOI2BB2X1 U785 ( .B0(N842), .B1(n638), .A0N(n634), .A1N(n746), .Y(n748) );
  AOI2BB2X1 U786 ( .B0(N481), .B1(n642), .A0N(n330), .A1N(n640), .Y(n747) );
  NAND2X1 U787 ( .A(n751), .B(n750), .Y(n457) );
  AOI2BB2X1 U788 ( .B0(N841), .B1(n638), .A0N(n634), .A1N(n749), .Y(n751) );
  AOI2BB2X1 U789 ( .B0(N480), .B1(n642), .A0N(n329), .A1N(n834), .Y(n750) );
  NAND2X1 U790 ( .A(n754), .B(n753), .Y(n458) );
  AOI2BB2X1 U791 ( .B0(N840), .B1(n638), .A0N(n635), .A1N(n752), .Y(n754) );
  AOI2BB2X1 U792 ( .B0(N479), .B1(n642), .A0N(n328), .A1N(n834), .Y(n753) );
  NAND2X1 U793 ( .A(n757), .B(n756), .Y(n459) );
  AOI2BB2X1 U794 ( .B0(N839), .B1(n638), .A0N(n635), .A1N(n755), .Y(n757) );
  AOI2BB2X1 U795 ( .B0(N478), .B1(n642), .A0N(n327), .A1N(n640), .Y(n756) );
  NAND2X1 U796 ( .A(n733), .B(n732), .Y(n451) );
  AOI2BB2X1 U797 ( .B0(N847), .B1(n638), .A0N(n634), .A1N(n731), .Y(n733) );
  AOI2BB2X1 U798 ( .B0(N486), .B1(n642), .A0N(n335), .A1N(n639), .Y(n732) );
  OAI211X1 U799 ( .A0(n661), .A1(n660), .B0(n869), .C0(n659), .Y(next_State[0]) );
  OA22X1 U800 ( .A0(n79), .A1(n686), .B0(n622), .B1(n704), .Y(n659) );
  OA22X1 U801 ( .A0(n423), .A1(n669), .B0(n244), .B1(n866), .Y(n661) );
  NOR2X1 U802 ( .A(ready), .B(n865), .Y(n244) );
  OAI222XL U803 ( .A0(index_X_After[0]), .A1(n869), .B0(n395), .B1(n623), .C0(
        n439), .C1(n628), .Y(n484) );
  OAI222XL U804 ( .A0(n395), .A1(n869), .B0(n394), .B1(n623), .C0(n438), .C1(
        n628), .Y(n485) );
  OAI222XL U805 ( .A0(n394), .A1(n869), .B0(n393), .B1(n623), .C0(n437), .C1(
        n628), .Y(n486) );
  OAI222XL U806 ( .A0(n393), .A1(n869), .B0(n392), .B1(n623), .C0(n436), .C1(
        n628), .Y(n487) );
  OAI222XL U807 ( .A0(n392), .A1(n869), .B0(n391), .B1(n623), .C0(n435), .C1(
        n628), .Y(n488) );
  OAI222XL U808 ( .A0(n391), .A1(n869), .B0(n401), .B1(n623), .C0(n434), .C1(
        n628), .Y(n489) );
  OAI222XL U809 ( .A0(n402), .A1(n869), .B0(n400), .B1(n623), .C0(n433), .C1(
        n628), .Y(n490) );
  OAI222XL U810 ( .A0(n401), .A1(n869), .B0(n399), .B1(n623), .C0(n432), .C1(
        n628), .Y(n491) );
  OAI222XL U811 ( .A0(n400), .A1(n869), .B0(n398), .B1(n623), .C0(n431), .C1(
        n628), .Y(n492) );
  OAI222XL U812 ( .A0(n399), .A1(n869), .B0(n397), .B1(n623), .C0(n430), .C1(
        n628), .Y(n493) );
  NAND2X1 U813 ( .A(n763), .B(n762), .Y(n461) );
  AOI2BB2X1 U814 ( .B0(N837), .B1(n637), .A0N(n635), .A1N(n761), .Y(n763) );
  AOI2BB2X1 U815 ( .B0(N476), .B1(n642), .A0N(n325), .A1N(n640), .Y(n762) );
  NAND2X1 U816 ( .A(n766), .B(n765), .Y(n462) );
  AOI2BB2X1 U817 ( .B0(N836), .B1(n637), .A0N(n635), .A1N(n764), .Y(n766) );
  AOI2BB2X1 U818 ( .B0(N475), .B1(n641), .A0N(n324), .A1N(n640), .Y(n765) );
  NAND2X1 U819 ( .A(n769), .B(n768), .Y(n463) );
  AOI2BB2X1 U820 ( .B0(N835), .B1(n637), .A0N(n635), .A1N(n767), .Y(n769) );
  AOI2BB2X1 U821 ( .B0(N474), .B1(n641), .A0N(n323), .A1N(n640), .Y(n768) );
  NAND2X1 U822 ( .A(n772), .B(n771), .Y(n464) );
  AOI2BB2X1 U823 ( .B0(N834), .B1(n637), .A0N(n635), .A1N(n770), .Y(n772) );
  AOI2BB2X1 U824 ( .B0(N473), .B1(n641), .A0N(n322), .A1N(n640), .Y(n771) );
  NAND2X1 U825 ( .A(n781), .B(n780), .Y(n467) );
  AOI2BB2X1 U826 ( .B0(N831), .B1(n637), .A0N(n635), .A1N(n779), .Y(n781) );
  AOI2BB2X1 U827 ( .B0(N470), .B1(n641), .A0N(n319), .A1N(n640), .Y(n780) );
  NAND2X1 U828 ( .A(n784), .B(n783), .Y(n468) );
  AOI2BB2X1 U829 ( .B0(N830), .B1(n637), .A0N(n635), .A1N(n782), .Y(n784) );
  AOI2BB2X1 U830 ( .B0(N469), .B1(n641), .A0N(n318), .A1N(n640), .Y(n783) );
  OAI22XL U831 ( .A0(n302), .A1(n628), .B0(n398), .B1(n869), .Y(n494) );
  OAI22XL U832 ( .A0(n301), .A1(n628), .B0(n397), .B1(n869), .Y(n495) );
  NAND2X1 U834 ( .A(n623), .B(n238), .Y(n508) );
  OAI21XL U835 ( .A0(n865), .A1(n424), .B0(n950), .Y(n238) );
  NAND3X1 U836 ( .A(n78), .B(n79), .C(n373), .Y(n388) );
  NAND3X1 U837 ( .A(n80), .B(n865), .C(next_State[0]), .Y(n78) );
  NAND2X1 U838 ( .A(n775), .B(n774), .Y(n465) );
  AOI2BB2X1 U839 ( .B0(N833), .B1(n637), .A0N(n635), .A1N(n773), .Y(n775) );
  AOI2BB2X1 U840 ( .B0(N472), .B1(n641), .A0N(n321), .A1N(n640), .Y(n774) );
  NAND2X1 U841 ( .A(n778), .B(n777), .Y(n466) );
  AOI2BB2X1 U842 ( .B0(N832), .B1(n637), .A0N(n635), .A1N(n776), .Y(n778) );
  AOI2BB2X1 U843 ( .B0(N471), .B1(n641), .A0N(n320), .A1N(n640), .Y(n777) );
  NAND2X1 U844 ( .A(n787), .B(n786), .Y(n469) );
  AOI2BB2X1 U845 ( .B0(N829), .B1(n637), .A0N(n635), .A1N(n785), .Y(n787) );
  AOI2BB2X1 U846 ( .B0(N468), .B1(n641), .A0N(n317), .A1N(n640), .Y(n786) );
  NAND2X1 U847 ( .A(n790), .B(n789), .Y(n470) );
  AOI2BB2X1 U848 ( .B0(N828), .B1(n637), .A0N(n636), .A1N(n788), .Y(n790) );
  AOI2BB2X1 U849 ( .B0(N467), .B1(n641), .A0N(n316), .A1N(n640), .Y(n789) );
  NAND2X1 U850 ( .A(n793), .B(n792), .Y(n471) );
  AOI2BB2X1 U851 ( .B0(N827), .B1(n637), .A0N(n636), .A1N(n791), .Y(n793) );
  AOI2BB2X1 U852 ( .B0(N466), .B1(n641), .A0N(n315), .A1N(n640), .Y(n792) );
  NAND2X1 U853 ( .A(n796), .B(n795), .Y(n472) );
  AOI2BB2X1 U854 ( .B0(N826), .B1(n613), .A0N(n636), .A1N(n794), .Y(n796) );
  AOI2BB2X1 U855 ( .B0(N465), .B1(n641), .A0N(n314), .A1N(n640), .Y(n795) );
  NAND2X1 U856 ( .A(n805), .B(n804), .Y(n475) );
  AOI2BB2X1 U857 ( .B0(N823), .B1(n613), .A0N(n636), .A1N(n803), .Y(n805) );
  AOI2BB2X1 U858 ( .B0(N462), .B1(n641), .A0N(n311), .A1N(n639), .Y(n804) );
  OAI21XL U859 ( .A0(n429), .A1(n247), .B0(n881), .Y(n510) );
  NOR3X1 U860 ( .A(n866), .B(n423), .C(n424), .Y(n247) );
  CLKINVX1 U861 ( .A(ready), .Y(n881) );
  NAND2X1 U862 ( .A(n799), .B(n798), .Y(n473) );
  AOI2BB2X1 U863 ( .B0(N825), .B1(n613), .A0N(n636), .A1N(n797), .Y(n799) );
  AOI2BB2X1 U864 ( .B0(N464), .B1(n642), .A0N(n313), .A1N(n639), .Y(n798) );
  NAND2X1 U865 ( .A(n802), .B(n801), .Y(n474) );
  AOI2BB2X1 U866 ( .B0(N824), .B1(n637), .A0N(n636), .A1N(n800), .Y(n802) );
  AOI2BB2X1 U867 ( .B0(N463), .B1(n530), .A0N(n312), .A1N(n639), .Y(n801) );
  NAND2X1 U868 ( .A(n808), .B(n807), .Y(n476) );
  AOI2BB2X1 U869 ( .B0(N822), .B1(n638), .A0N(n636), .A1N(n806), .Y(n808) );
  AOI2BB2X1 U870 ( .B0(N461), .B1(n530), .A0N(n310), .A1N(n639), .Y(n807) );
  NAND2X1 U871 ( .A(n811), .B(n810), .Y(n477) );
  AOI2BB2X1 U872 ( .B0(N821), .B1(n637), .A0N(n636), .A1N(n809), .Y(n811) );
  AOI2BB2X1 U873 ( .B0(N460), .B1(n530), .A0N(n309), .A1N(n639), .Y(n810) );
  NAND2X1 U874 ( .A(n814), .B(n813), .Y(n478) );
  AOI2BB2X1 U875 ( .B0(N820), .B1(n638), .A0N(n636), .A1N(n812), .Y(n814) );
  AOI2BB2X1 U876 ( .B0(N459), .B1(n530), .A0N(n308), .A1N(n639), .Y(n813) );
  NAND2X1 U877 ( .A(n820), .B(n819), .Y(n480) );
  AOI2BB2X1 U878 ( .B0(N818), .B1(n637), .A0N(n636), .A1N(n818), .Y(n820) );
  AOI2BB2X1 U879 ( .B0(N457), .B1(n530), .A0N(n306), .A1N(n639), .Y(n819) );
  NAND2X1 U880 ( .A(n826), .B(n825), .Y(n482) );
  AOI2BB2X1 U881 ( .B0(N455), .B1(n530), .A0N(n304), .A1N(n639), .Y(n825) );
  AOI2BB2X1 U882 ( .B0(N816), .B1(n638), .A0N(n635), .A1N(n824), .Y(n826) );
  NAND2X1 U883 ( .A(n829), .B(n828), .Y(n483) );
  AOI2BB2X1 U884 ( .B0(N454), .B1(n530), .A0N(n303), .A1N(n639), .Y(n828) );
  AOI2BB2X1 U885 ( .B0(N815), .B1(n637), .A0N(n636), .A1N(n827), .Y(n829) );
  NAND2X1 U886 ( .A(n817), .B(n816), .Y(n479) );
  AOI2BB2X1 U887 ( .B0(N819), .B1(n638), .A0N(n636), .A1N(n815), .Y(n817) );
  AOI2BB2X1 U888 ( .B0(N458), .B1(n530), .A0N(n307), .A1N(n639), .Y(n816) );
  NAND2X1 U889 ( .A(n823), .B(n822), .Y(n481) );
  AOI2BB2X1 U890 ( .B0(N456), .B1(n530), .A0N(n305), .A1N(n639), .Y(n822) );
  AOI2BB2X1 U891 ( .B0(N817), .B1(n637), .A0N(n636), .A1N(n821), .Y(n823) );
  OAI22XL U892 ( .A0(n370), .A1(n624), .B0(n43), .B1(n622), .Y(n379) );
  AOI222XL U893 ( .A0(index_X_After[3]), .A1(n843), .B0(index_X[3]), .B1(n842), 
        .C0(index_X_Before[3]), .C1(n841), .Y(n43) );
  NAND2X1 U894 ( .A(n423), .B(n660), .Y(n79) );
  OAI22XL U895 ( .A0(n371), .A1(n624), .B0(n45), .B1(n622), .Y(n380) );
  AOI222XL U896 ( .A0(index_X_After[4]), .A1(n843), .B0(n890), .B1(n842), .C0(
        index_X_Before[4]), .C1(n841), .Y(n45) );
  NAND3BX1 U897 ( .AN(n374), .B(n423), .C(n662), .Y(n668) );
  OAI221XL U898 ( .A0(n895), .A1(n864), .B0(n624), .B1(n592), .C0(n859), .Y(
        n385) );
  AOI2BB2X1 U899 ( .B0(index_Y_Before[3]), .B1(n862), .A0N(n399), .A1N(n861), 
        .Y(n859) );
  OAI221XL U900 ( .A0(n892), .A1(n864), .B0(n624), .B1(n576), .C0(n863), .Y(
        n387) );
  AOI2BB2X1 U901 ( .B0(index_Y_Before[5]), .B1(n862), .A0N(n397), .A1N(n861), 
        .Y(n863) );
  NAND4X1 U902 ( .A(n392), .B(n393), .C(n391), .D(n224), .Y(n210) );
  NOR3X1 U903 ( .A(n891), .B(N144), .C(n889), .Y(n224) );
  OAI22XL U904 ( .A0(n372), .A1(n624), .B0(n47), .B1(n622), .Y(n381) );
  AOI222XL U905 ( .A0(index_X_After[5]), .A1(n843), .B0(index_X[5]), .B1(n842), 
        .C0(index_X_Before[5]), .C1(n841), .Y(n47) );
  OAI22XL U906 ( .A0(n367), .A1(n624), .B0(n34), .B1(n622), .Y(n376) );
  AOI222XL U907 ( .A0(index_X_After[0]), .A1(n843), .B0(N144), .B1(n842), .C0(
        index_X_After[0]), .C1(n841), .Y(n34) );
  OAI22XL U908 ( .A0(n368), .A1(n624), .B0(n39), .B1(n622), .Y(n377) );
  AOI222XL U909 ( .A0(index_X_After[1]), .A1(n843), .B0(n889), .B1(n842), .C0(
        index_X_Before[1]), .C1(n841), .Y(n39) );
  OAI22XL U910 ( .A0(n369), .A1(n624), .B0(n41), .B1(n622), .Y(n378) );
  AOI222XL U911 ( .A0(index_X_After[2]), .A1(n843), .B0(n891), .B1(n842), .C0(
        index_X_Before[2]), .C1(n841), .Y(n41) );
  NOR4X1 U912 ( .A(n220), .B(index_Y[5]), .C(index_Y[3]), .D(n893), .Y(n213)
         );
  NAND3X1 U913 ( .A(n401), .B(n402), .C(n400), .Y(n220) );
  NOR2BX1 U914 ( .AN(n219), .B(n402), .Y(n30) );
  CLKBUFX3 U915 ( .A(n24), .Y(n622) );
  NAND3BX1 U916 ( .AN(n865), .B(n424), .C(n866), .Y(n24) );
  OAI21XL U917 ( .A0(n399), .A1(n257), .B0(n261), .Y(n517) );
  AOI22X1 U918 ( .A0(N178), .A1(n259), .B0(n260), .B1(index_Y_After[3]), .Y(
        n261) );
  OAI21XL U919 ( .A0(n400), .A1(n257), .B0(n262), .Y(n518) );
  AOI22X1 U920 ( .A0(N177), .A1(n259), .B0(n260), .B1(index_Y_After[2]), .Y(
        n262) );
  OAI21XL U921 ( .A0(n401), .A1(n257), .B0(n263), .Y(n519) );
  AOI22X1 U922 ( .A0(N176), .A1(n259), .B0(n260), .B1(index_Y_After[1]), .Y(
        n263) );
  CLKINVX1 U923 ( .A(index_Y[1]), .Y(N176) );
  OAI21XL U924 ( .A0(n402), .A1(n257), .B0(n264), .Y(n520) );
  AOI22X1 U925 ( .A0(N175), .A1(n259), .B0(n260), .B1(n402), .Y(n264) );
  OAI21XL U926 ( .A0(n398), .A1(n257), .B0(n258), .Y(n516) );
  AOI22X1 U927 ( .A0(N179), .A1(n259), .B0(n260), .B1(index_Y_After[4]), .Y(
        n258) );
  OAI21XL U928 ( .A0(n397), .A1(n257), .B0(n267), .Y(n522) );
  AOI22X1 U929 ( .A0(N180), .A1(n259), .B0(n260), .B1(index_Y_After[5]), .Y(
        n267) );
  AND4X1 U930 ( .A(n890), .B(index_X[5]), .C(index_X[3]), .D(n269), .Y(n268)
         );
  NOR2X1 U931 ( .A(n394), .B(n395), .Y(n269) );
  CLKINVX1 U932 ( .A(n394), .Y(n891) );
  CLKINVX1 U933 ( .A(n395), .Y(n889) );
  CLKINVX1 U934 ( .A(n398), .Y(n893) );
  AND4X1 U935 ( .A(n893), .B(index_Y[5]), .C(index_Y[3]), .D(n246), .Y(n219)
         );
  NOR2X1 U936 ( .A(n400), .B(n401), .Y(n246) );
  CLKINVX1 U937 ( .A(n392), .Y(n890) );
  NAND2X1 U938 ( .A(n620), .B(n604), .Y(n845) );
  NAND2X1 U939 ( .A(n620), .B(n609), .Y(n847) );
  OAI222XL U940 ( .A0(index_X_After[0]), .A1(n845), .B0(N144), .B1(n844), .C0(
        n300), .C1(n627), .Y(n496) );
  OAI222XL U941 ( .A0(n395), .A1(n845), .B0(n888), .B1(n844), .C0(n299), .C1(
        n627), .Y(n497) );
  OAI222XL U942 ( .A0(n394), .A1(n845), .B0(n887), .B1(n844), .C0(n298), .C1(
        n627), .Y(n498) );
  OAI222XL U943 ( .A0(n393), .A1(n845), .B0(n886), .B1(n844), .C0(n297), .C1(
        n627), .Y(n499) );
  OAI222XL U944 ( .A0(n392), .A1(n845), .B0(n885), .B1(n844), .C0(n296), .C1(
        n627), .Y(n500) );
  OAI222XL U945 ( .A0(n391), .A1(n845), .B0(n884), .B1(n844), .C0(n295), .C1(
        n627), .Y(n501) );
  OAI222XL U946 ( .A0(n402), .A1(n847), .B0(N175), .B1(n846), .C0(n294), .C1(
        n627), .Y(n502) );
  OAI222XL U947 ( .A0(n401), .A1(n847), .B0(n897), .B1(n846), .C0(n293), .C1(
        n627), .Y(n503) );
  OAI222XL U948 ( .A0(n400), .A1(n847), .B0(n896), .B1(n846), .C0(n292), .C1(
        n627), .Y(n504) );
  OAI222XL U949 ( .A0(n399), .A1(n847), .B0(n895), .B1(n846), .C0(n291), .C1(
        n627), .Y(n505) );
  OAI222XL U950 ( .A0(n398), .A1(n847), .B0(n894), .B1(n846), .C0(n290), .C1(
        n627), .Y(n506) );
  OAI222XL U951 ( .A0(n397), .A1(n847), .B0(n892), .B1(n846), .C0(n289), .C1(
        n627), .Y(n507) );
  OAI221XL U952 ( .A0(n897), .A1(n864), .B0(n624), .B1(n582), .C0(n857), .Y(
        n383) );
  AOI2BB2X1 U953 ( .B0(index_Y_Before[1]), .B1(n862), .A0N(n401), .A1N(n861), 
        .Y(n857) );
  OAI221XL U954 ( .A0(n896), .A1(n864), .B0(n624), .B1(n580), .C0(n858), .Y(
        n384) );
  AOI2BB2X1 U955 ( .B0(index_Y_Before[2]), .B1(n862), .A0N(n400), .A1N(n861), 
        .Y(n858) );
  OAI221XL U956 ( .A0(n894), .A1(n864), .B0(n624), .B1(n578), .C0(n860), .Y(
        n386) );
  AOI2BB2X1 U957 ( .B0(index_Y_Before[4]), .B1(n862), .A0N(n398), .A1N(n861), 
        .Y(n860) );
  OAI221XL U958 ( .A0(n870), .A1(n686), .B0(n622), .B1(n690), .C0(n658), .Y(
        next_State[1]) );
  AOI31X1 U959 ( .A0(n26), .A1(n374), .A2(n660), .B0(n657), .Y(n658) );
  CLKINVX1 U960 ( .A(n29), .Y(n657) );
  AO21X1 U961 ( .A0(n30), .A1(n883), .B0(n865), .Y(n26) );
  OAI221XL U962 ( .A0(n670), .A1(n668), .B0(n609), .B1(n667), .C0(n674), .Y(
        n524) );
  OAI221XL U963 ( .A0(n886), .A1(n249), .B0(n393), .B1(n250), .C0(n253), .Y(
        n512) );
  NAND2X1 U964 ( .A(N147), .B(n252), .Y(n253) );
  OAI221XL U965 ( .A0(n887), .A1(n249), .B0(n394), .B1(n250), .C0(n254), .Y(
        n513) );
  NAND2X1 U966 ( .A(N146), .B(n252), .Y(n254) );
  OAI221XL U967 ( .A0(n885), .A1(n249), .B0(n392), .B1(n250), .C0(n251), .Y(
        n511) );
  NAND2X1 U968 ( .A(N148), .B(n252), .Y(n251) );
  OAI221XL U969 ( .A0(n888), .A1(n249), .B0(n395), .B1(n250), .C0(n255), .Y(
        n514) );
  NAND2X1 U970 ( .A(N145), .B(n252), .Y(n255) );
  CLKINVX1 U971 ( .A(index_X[1]), .Y(N145) );
  OAI221XL U972 ( .A0(N144), .A1(n249), .B0(index_X_After[0]), .B1(n250), .C0(
        n256), .Y(n515) );
  NAND2X1 U973 ( .A(N144), .B(n252), .Y(n256) );
  OAI221XL U974 ( .A0(n884), .A1(n249), .B0(n391), .B1(n250), .C0(n265), .Y(
        n521) );
  NAND2X1 U975 ( .A(N149), .B(n252), .Y(n265) );
  OAI221XL U976 ( .A0(n856), .A1(N175), .B0(n402), .B1(n861), .C0(n855), .Y(
        n382) );
  OA22X1 U977 ( .A0(N175), .A1(n864), .B0(n624), .B1(n584), .Y(n855) );
  NAND2X1 U978 ( .A(index_X_After[0]), .B(n268), .Y(n245) );
  AO21X1 U979 ( .A0(n424), .A1(n669), .B0(n374), .Y(n80) );
  AND2X2 U980 ( .A(n346), .B(n266), .Y(n621) );
  NOR2X1 U981 ( .A(n79), .B(n374), .Y(n229) );
  CLKINVX1 U982 ( .A(n239), .Y(n669) );
  NAND3BX1 U983 ( .AN(n245), .B(n219), .C(n402), .Y(n239) );
  CLKINVX1 U984 ( .A(index_X[3]), .Y(n875) );
  CLKINVX1 U985 ( .A(index_Y[3]), .Y(n880) );
  NAND2X1 U986 ( .A(n375), .B(n870), .Y(n389) );
  OR2X4 U987 ( .A(n671), .B(N363), .Y(n104) );
  XOR2X1 U988 ( .A(index_Y[5]), .B(\add_112_S2/carry[5] ), .Y(N180) );
  AND2X1 U989 ( .A(\add_112_S2/carry[4] ), .B(index_Y[4]), .Y(
        \add_112_S2/carry[5] ) );
  XOR2X1 U990 ( .A(index_Y[4]), .B(\add_112_S2/carry[4] ), .Y(N179) );
  AND2X1 U991 ( .A(\add_112_S2/carry[3] ), .B(index_Y[3]), .Y(
        \add_112_S2/carry[4] ) );
  XOR2X1 U992 ( .A(index_Y[3]), .B(\add_112_S2/carry[3] ), .Y(N178) );
  AND2X1 U993 ( .A(index_Y[1]), .B(index_Y[2]), .Y(\add_112_S2/carry[3] ) );
  XOR2X1 U994 ( .A(index_Y[2]), .B(index_Y[1]), .Y(N177) );
  XOR2X1 U995 ( .A(index_X[5]), .B(\add_99/carry[5] ), .Y(N149) );
  AND2X1 U996 ( .A(\add_99/carry[4] ), .B(index_X[4]), .Y(\add_99/carry[5] )
         );
  XOR2X1 U997 ( .A(index_X[4]), .B(\add_99/carry[4] ), .Y(N148) );
  AND2X1 U998 ( .A(\add_99/carry[3] ), .B(index_X[3]), .Y(\add_99/carry[4] )
         );
  XOR2X1 U999 ( .A(index_X[3]), .B(\add_99/carry[3] ), .Y(N147) );
  AND2X1 U1000 ( .A(index_X[1]), .B(index_X[2]), .Y(\add_99/carry[3] ) );
  XOR2X1 U1001 ( .A(index_X[2]), .B(index_X[1]), .Y(N146) );
  XOR2X1 U1002 ( .A(\r354/carry[5] ), .B(index_X[5]), .Y(index_X_After[5]) );
  XOR2X1 U1003 ( .A(\r356/carry[5] ), .B(index_Y[5]), .Y(index_Y_After[5]) );
  NAND2BX1 U1004 ( .AN(index_X[1]), .B(index_X_After[0]), .Y(n871) );
  OAI2BB1X1 U1005 ( .A0N(N144), .A1N(index_X[1]), .B0(n871), .Y(
        index_X_Before[1]) );
  NOR2X1 U1006 ( .A(n871), .B(index_X[2]), .Y(n872) );
  AO21X1 U1007 ( .A0(n871), .A1(index_X[2]), .B0(n872), .Y(index_X_Before[2])
         );
  NAND2X1 U1008 ( .A(n872), .B(n875), .Y(n873) );
  OAI21XL U1009 ( .A0(n872), .A1(n875), .B0(n873), .Y(index_X_Before[3]) );
  XNOR2X1 U1010 ( .A(index_X[4]), .B(n873), .Y(index_X_Before[4]) );
  NOR2X1 U1011 ( .A(index_X[4]), .B(n873), .Y(n874) );
  XOR2X1 U1012 ( .A(index_X[5]), .B(n874), .Y(index_X_Before[5]) );
  NAND2BX1 U1013 ( .AN(index_Y[1]), .B(n402), .Y(n876) );
  OAI2BB1X1 U1014 ( .A0N(N175), .A1N(index_Y[1]), .B0(n876), .Y(
        index_Y_Before[1]) );
  NOR2X1 U1015 ( .A(n876), .B(index_Y[2]), .Y(n877) );
  AO21X1 U1016 ( .A0(n876), .A1(index_Y[2]), .B0(n877), .Y(index_Y_Before[2])
         );
  NAND2X1 U1017 ( .A(n877), .B(n880), .Y(n878) );
  OAI21XL U1018 ( .A0(n877), .A1(n880), .B0(n878), .Y(index_Y_Before[3]) );
  XNOR2X1 U1019 ( .A(index_Y[4]), .B(n878), .Y(index_Y_Before[4]) );
  NOR2X1 U1020 ( .A(index_Y[4]), .B(n878), .Y(n879) );
  XOR2X1 U1021 ( .A(index_Y[5]), .B(n879), .Y(index_Y_Before[5]) );
  CONV_DW01_add_0 add_286 ( .A(convTemp), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N858, N857, N856, N855, N854, 
        N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, 
        N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, 
        N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, 
        N817, N816, N815}) );
  CONV_DW_cmp_0 gt_259 ( .A(cdata_rd), .B({n917, cdata_wr[18], n919, n920, 
        cdata_wr[15], n922, cdata_wr[13], n924, cdata_wr[11], n926, 
        cdata_wr[9], n928, n929, cdata_wr[6], n931, cdata_wr[4], n933, n934, 
        cdata_wr[1:0]}), .TC(1'b0), .GE_LT(1'b0), .GE_GT_EQ(1'b1), 
        .GE_LT_GT_LE(N363) );
  CONV_DW01_inc_0 add_38 ( .A(convTemp[35:15]), .SUM({roundTemp, 
        SYNOPSYS_UNCONNECTED__0}) );
  CONV_DW_mult_tc_2 mult_266 ( .a({N53, N53, N53, N53, N61, N71, N78, N85, N89, 
        N90, N94, n882, N98, N102, N109, N111, N55, N114, N124, N128}), .b(
        idataTemp), .product({mulTemp_43, mulTemp}) );
  CONV_DW01_add_5 r362 ( .A(convTemp), .B({mulTemp_43, mulTemp_43, mulTemp_43, 
        mulTemp_43, mulTemp_43, mulTemp[38:16], n534, mulTemp[14:7], n527, 
        mulTemp[5:0]}), .CI(1'b0), .SUM({N497, N496, N495, N494, N493, N492, 
        N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, 
        N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, 
        N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, 
        N455, N454}) );
  DFFRXL \iaddr_reg[6]  ( .D(n382), .CK(clk), .RN(n868), .Q(n971), .QN(n584)
         );
  DFFRXL \iaddr_reg[11]  ( .D(n387), .CK(clk), .RN(n868), .Q(n966), .QN(n576)
         );
  DFFRXL \iaddr_reg[10]  ( .D(n386), .CK(clk), .RN(n868), .Q(n967), .QN(n578)
         );
  DFFRXL \iaddr_reg[9]  ( .D(n385), .CK(clk), .RN(n868), .Q(n968), .QN(n592)
         );
  DFFRXL \iaddr_reg[8]  ( .D(n384), .CK(clk), .RN(n868), .Q(n969), .QN(n580)
         );
  DFFRXL \iaddr_reg[7]  ( .D(n383), .CK(clk), .RN(n868), .Q(n970), .QN(n582)
         );
  DFFRXL cwr_reg ( .D(n509), .CK(clk), .RN(n868), .Q(n972) );
  DFFRX2 \index_X_reg[0]  ( .D(n515), .CK(clk), .RN(n868), .Q(N144), .QN(
        index_X_After[0]) );
  INVX3 U490 ( .A(reset), .Y(n868) );
  INVXL U491 ( .A(n972), .Y(n952) );
  INVX12 U542 ( .A(n952), .Y(cwr) );
  INVXL U543 ( .A(n970), .Y(n954) );
  INVX12 U544 ( .A(n954), .Y(iaddr[7]) );
  INVXL U545 ( .A(n969), .Y(n956) );
  INVX12 U546 ( .A(n956), .Y(iaddr[8]) );
  INVXL U553 ( .A(n968), .Y(n958) );
  INVX12 U833 ( .A(n958), .Y(iaddr[9]) );
  INVXL U1022 ( .A(n967), .Y(n960) );
  INVX12 U1023 ( .A(n960), .Y(iaddr[10]) );
  INVXL U1024 ( .A(n966), .Y(n962) );
  INVX12 U1025 ( .A(n962), .Y(iaddr[11]) );
  INVXL U1026 ( .A(n971), .Y(n964) );
  INVX12 U1027 ( .A(n964), .Y(iaddr[6]) );
endmodule

